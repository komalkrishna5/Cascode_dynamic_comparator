magic
tech sky130A
timestamp 1654337383
<< error_s >>
rect 297 2301 326 2401
rect 341 2301 370 2401
rect 495 2302 524 2402
rect 539 2302 568 2402
rect 145 1373 174 1473
rect 189 1373 218 1473
rect 698 1373 727 1473
rect 742 1373 771 1473
<< nwell >>
rect 391 2526 470 2668
rect -57 1756 74 1784
rect -57 1574 843 1756
rect -57 1565 64 1574
rect 32 1178 159 1179
rect 32 1177 328 1178
rect 32 1152 179 1177
rect 220 1152 328 1177
rect 32 997 328 1152
rect 32 990 196 997
rect 32 966 167 990
rect 32 961 196 966
rect 232 961 328 997
rect 610 1004 658 1023
rect 610 996 655 1004
rect 32 840 328 961
rect 555 982 655 996
rect 555 980 658 982
rect 555 951 570 980
rect 610 967 658 980
rect 32 828 132 840
rect 195 831 328 840
rect 195 828 223 831
rect 32 808 353 828
rect 367 287 433 413
<< psubdiff >>
rect 43 -499 79 -487
rect 43 -575 79 -563
<< nsubdiff >>
rect 405 2635 444 2647
rect 405 2533 444 2545
rect -21 1712 13 1724
rect -21 1638 13 1650
rect 63 1144 122 1156
rect 63 1032 122 1044
rect 379 391 413 403
rect 379 317 413 329
<< psubdiffcont >>
rect 43 -563 79 -499
<< nsubdiffcont >>
rect 405 2545 444 2635
rect -21 1650 13 1712
rect 63 1044 122 1144
rect 379 329 413 391
<< poly >>
rect 326 2406 341 2410
rect 183 2303 221 2315
rect 183 2279 192 2303
rect 213 2289 221 2303
rect 684 2290 721 2300
rect 684 2289 692 2290
rect 213 2279 341 2289
rect 183 2266 341 2279
rect 524 2266 692 2289
rect 713 2266 721 2290
rect 684 2259 721 2266
rect 380 1934 492 1945
rect 380 1899 414 1934
rect 464 1899 492 1934
rect 380 1739 492 1899
rect 861 1608 896 1615
rect 783 1605 896 1608
rect 783 1588 870 1605
rect 887 1588 896 1605
rect 861 1578 896 1588
rect 174 1351 189 1366
rect 727 1355 742 1367
rect 618 1001 654 1012
rect 190 986 226 997
rect 618 996 626 1001
rect 190 969 198 986
rect 216 985 226 986
rect 216 969 279 985
rect 190 961 226 969
rect 264 933 279 969
rect 555 984 626 996
rect 644 984 654 1001
rect 555 980 654 984
rect 555 951 570 980
rect 618 976 654 980
rect 154 783 169 838
rect 264 831 279 832
rect 555 828 570 831
rect 664 790 679 830
rect 133 767 194 783
rect 133 744 150 767
rect 175 744 194 767
rect 133 729 194 744
rect 641 769 702 790
rect 641 744 657 769
rect 685 744 702 769
rect 641 736 702 744
rect 34 225 104 248
rect 34 202 53 225
rect 85 202 104 225
rect 748 225 818 248
rect 748 223 767 225
rect 34 180 104 202
rect 735 202 767 223
rect 799 202 818 225
rect 735 199 818 202
rect 748 180 818 199
<< polycont >>
rect 192 2279 213 2303
rect 692 2266 713 2290
rect 414 1899 464 1934
rect 870 1588 887 1605
rect 198 969 216 986
rect 626 984 644 1001
rect 150 744 175 767
rect 657 744 685 769
rect 53 202 85 225
rect 767 202 799 225
<< locali >>
rect -1296 2676 -675 2757
rect 1594 2727 2192 2778
rect 1594 2707 1640 2727
rect 1593 2705 1640 2707
rect 1306 2704 1640 2705
rect 198 2699 1640 2704
rect -1296 2319 -673 2676
rect 411 2643 440 2687
rect 574 2676 1640 2699
rect 405 2635 444 2643
rect 405 2537 444 2545
rect 1594 2607 1640 2676
rect 1752 2607 2040 2727
rect 2152 2607 2192 2727
rect 1594 2505 2192 2607
rect 257 2426 388 2460
rect 545 2431 595 2468
rect -1296 2146 -1256 2319
rect -1131 2146 -856 2319
rect -731 2254 -673 2319
rect 184 2305 221 2313
rect 184 2277 190 2305
rect 215 2277 221 2305
rect 184 2272 221 2277
rect 684 2291 721 2300
rect 684 2265 691 2291
rect 714 2265 721 2291
rect 684 2259 721 2265
rect -731 2227 212 2254
rect -731 2146 -673 2227
rect -1296 2045 -673 2146
rect -1296 1948 -681 2045
rect -1296 1413 -673 1948
rect 399 1934 477 1946
rect 399 1899 414 1934
rect 464 1899 477 1934
rect 399 1889 477 1899
rect -25 1849 16 1855
rect -25 1819 -19 1849
rect 10 1819 16 1849
rect -25 1811 16 1819
rect 1587 1848 2192 2505
rect -14 1720 5 1811
rect 1587 1728 1640 1848
rect 1752 1728 2040 1848
rect 2152 1728 2192 1848
rect -21 1712 13 1720
rect -21 1642 13 1650
rect 862 1608 895 1613
rect 862 1585 866 1608
rect 890 1585 895 1608
rect 862 1580 895 1585
rect -1296 1240 -1256 1413
rect -1131 1240 -856 1413
rect -731 1382 -673 1413
rect -731 1381 -17 1382
rect -731 1355 69 1381
rect -731 1240 -673 1355
rect -616 1354 -185 1355
rect 44 1344 69 1355
rect 44 1334 73 1344
rect -1296 -349 -673 1240
rect 1587 1242 2192 1728
rect 1587 1206 1640 1242
rect 1567 1205 1640 1206
rect 704 1204 927 1205
rect 1049 1204 1640 1205
rect 172 1193 218 1204
rect 127 1177 218 1193
rect 127 1152 179 1177
rect 63 1144 179 1152
rect -419 1009 -280 1057
rect 122 1055 179 1144
rect 122 1044 148 1055
rect 63 1036 148 1044
rect -419 964 -368 1009
rect -322 1000 -280 1009
rect -419 958 -322 964
rect -419 919 -280 958
rect 131 929 148 1036
rect 633 1015 655 1016
rect 610 1005 655 1015
rect 193 991 224 1000
rect 221 964 224 991
rect 610 980 620 1005
rect 648 980 655 1005
rect 610 973 655 980
rect 633 972 655 973
rect 193 958 224 964
rect 685 919 702 1189
rect 704 1178 1640 1204
rect 704 1177 1564 1178
rect 927 1176 1029 1177
rect 1587 1122 1640 1178
rect 1752 1122 2040 1242
rect 2152 1122 2192 1242
rect 1181 1016 1319 1057
rect 1232 1009 1319 1016
rect 1181 964 1232 972
rect 1278 964 1319 1009
rect 1181 919 1319 964
rect 133 770 194 783
rect 133 741 147 770
rect 178 741 194 770
rect 133 729 194 741
rect 641 776 702 790
rect 641 739 650 776
rect 695 739 702 776
rect 641 736 658 739
rect 681 736 702 739
rect 1587 716 2192 1122
rect 1587 543 2194 716
rect 825 462 1087 463
rect 1587 462 1640 543
rect 386 399 405 452
rect 825 434 1640 462
rect 1411 433 1640 434
rect 379 391 413 399
rect 1587 371 1640 433
rect 1752 371 2040 543
rect 2152 371 2194 543
rect 379 321 413 329
rect -406 291 -294 312
rect 1160 308 1335 333
rect -440 266 -265 291
rect -440 147 -407 266
rect -294 147 -265 266
rect 34 227 104 248
rect 34 200 51 227
rect 87 200 104 227
rect 34 180 104 200
rect 748 227 818 248
rect 748 200 765 227
rect 801 200 818 227
rect 748 180 818 200
rect 1160 199 1193 308
rect 1159 177 1193 199
rect 1306 177 1335 308
rect 1587 180 2194 371
rect 1159 170 1335 177
rect 1160 152 1335 170
rect -406 146 -294 147
rect 1589 83 2194 180
rect -1296 -522 -1256 -349
rect -1131 -522 -856 -349
rect -731 -443 -673 -349
rect -731 -444 -508 -443
rect -731 -469 13 -444
rect 60 -462 79 -448
rect -731 -522 -673 -469
rect -508 -470 13 -469
rect -1296 -765 -673 -522
rect 43 -499 79 -462
rect 43 -571 79 -563
rect -440 -614 -265 -589
rect -440 -745 -407 -614
rect -294 -638 -265 -614
rect 1590 -629 2192 83
rect -294 -745 -265 -724
rect -1296 -967 -675 -765
rect -440 -771 -265 -745
rect 1590 -965 2193 -629
<< viali >>
rect 1640 2607 1752 2727
rect 2040 2607 2152 2727
rect -1256 2146 -1131 2319
rect -856 2146 -731 2319
rect 190 2303 215 2305
rect 190 2279 192 2303
rect 192 2279 213 2303
rect 213 2279 215 2303
rect 190 2277 215 2279
rect 691 2290 714 2291
rect 691 2266 692 2290
rect 692 2266 713 2290
rect 713 2266 714 2290
rect 691 2265 714 2266
rect 414 1899 464 1934
rect -19 1819 10 1849
rect 1640 1728 1752 1848
rect 2040 1728 2152 1848
rect 866 1605 890 1608
rect 866 1588 870 1605
rect 870 1588 887 1605
rect 887 1588 890 1605
rect 866 1585 890 1588
rect -1256 1240 -1131 1413
rect -856 1240 -731 1413
rect -368 964 -322 1009
rect 193 986 221 991
rect 193 969 198 986
rect 198 969 216 986
rect 216 969 221 986
rect 193 964 221 969
rect 620 1001 648 1005
rect 620 984 626 1001
rect 626 984 644 1001
rect 644 984 648 1001
rect 620 980 648 984
rect 1640 1122 1752 1242
rect 2040 1122 2152 1242
rect 1232 964 1278 1009
rect 147 767 178 770
rect 147 744 150 767
rect 150 744 175 767
rect 175 744 178 767
rect 147 741 178 744
rect 650 769 695 776
rect 650 744 657 769
rect 657 744 685 769
rect 685 744 695 769
rect 650 739 695 744
rect 1640 371 1752 543
rect 2040 371 2152 543
rect -407 147 -294 266
rect 51 225 87 227
rect 51 202 53 225
rect 53 202 85 225
rect 85 202 87 225
rect 51 200 87 202
rect 765 225 801 227
rect 765 202 767 225
rect 767 202 799 225
rect 799 202 801 225
rect 765 200 801 202
rect 1193 177 1306 308
rect -1256 -522 -1131 -349
rect -856 -522 -731 -349
rect -407 -745 -294 -614
<< metal1 >>
rect 1605 2727 1783 2757
rect 1605 2607 1640 2727
rect 1752 2607 1783 2727
rect 1605 2574 1783 2607
rect 2004 2727 2183 2757
rect 2004 2607 2040 2727
rect 2152 2607 2183 2727
rect 2004 2574 2183 2607
rect -1285 2319 -1102 2342
rect -1285 2146 -1256 2319
rect -1131 2146 -1102 2319
rect -1285 2113 -1102 2146
rect -885 2319 -702 2342
rect -885 2146 -856 2319
rect -731 2146 -702 2319
rect 182 2305 222 2314
rect -885 2113 -702 2146
rect -159 2277 190 2305
rect 215 2277 222 2305
rect -159 1570 -119 2277
rect 182 2271 222 2277
rect 684 2291 721 2300
rect 684 2265 691 2291
rect 714 2290 721 2291
rect 714 2267 1029 2290
rect 714 2265 721 2267
rect 684 2259 721 2265
rect 381 2076 509 2111
rect 380 2014 412 2076
rect 480 2014 509 2076
rect 380 1984 509 2014
rect 380 1934 492 1984
rect 988 1961 1029 2267
rect 380 1899 414 1934
rect 464 1899 492 1934
rect 380 1886 492 1899
rect -25 1849 16 1855
rect 402 1851 521 1864
rect 402 1849 433 1851
rect -25 1819 -19 1849
rect 10 1819 433 1849
rect -25 1818 433 1819
rect -25 1811 16 1818
rect 402 1811 433 1818
rect 485 1811 521 1851
rect 402 1800 521 1811
rect 989 1616 1029 1961
rect 1604 1848 1783 1878
rect 1604 1728 1640 1848
rect 1752 1728 1783 1848
rect 1604 1695 1783 1728
rect 2004 1848 2183 1878
rect 2004 1728 2040 1848
rect 2152 1728 2183 1848
rect 2004 1695 2183 1728
rect 857 1608 1029 1616
rect 857 1585 866 1608
rect 890 1603 1029 1608
rect 890 1585 1031 1603
rect 857 1578 1031 1585
rect -159 1537 180 1570
rect -1285 1413 -1102 1438
rect -1285 1240 -1256 1413
rect -1131 1240 -1102 1413
rect -1285 1207 -1102 1240
rect -885 1413 -702 1438
rect -885 1240 -856 1413
rect -731 1240 -702 1413
rect -885 1207 -702 1240
rect -423 1018 -279 1056
rect -423 958 -375 1018
rect -315 958 -279 1018
rect -423 919 -279 958
rect -453 291 -266 311
rect -453 266 -265 291
rect -453 147 -407 266
rect -294 147 -265 266
rect -453 124 -266 147
rect -1285 -349 -1102 -324
rect -1285 -522 -1256 -349
rect -1131 -522 -1102 -349
rect -1285 -555 -1102 -522
rect -885 -349 -702 -324
rect -885 -522 -856 -349
rect -731 -522 -702 -349
rect -159 -368 -119 1537
rect 988 1300 1031 1578
rect 610 1007 655 1016
rect 187 991 227 1000
rect 187 964 193 991
rect 221 964 227 991
rect 610 978 619 1007
rect 650 978 655 1007
rect 610 973 655 978
rect 187 958 227 964
rect 133 773 194 783
rect 133 739 145 773
rect 180 739 194 773
rect 133 729 194 739
rect 283 691 303 890
rect -29 660 303 691
rect 528 697 552 867
rect 641 776 702 790
rect 641 739 650 776
rect 695 739 702 776
rect 641 736 702 739
rect -29 -290 -1 660
rect 528 658 941 697
rect 682 300 711 390
rect 34 230 104 248
rect 34 197 48 230
rect 90 197 104 230
rect 34 180 104 197
rect 682 118 707 300
rect 893 248 941 658
rect 988 313 1032 1300
rect 1604 1242 1783 1272
rect 1604 1122 1640 1242
rect 1752 1122 1783 1242
rect 1604 1091 1783 1122
rect 2004 1242 2183 1272
rect 2004 1122 2040 1242
rect 2152 1122 2183 1242
rect 2004 1091 2183 1122
rect 1177 1018 1319 1056
rect 1177 958 1225 1018
rect 1285 958 1319 1018
rect 1177 919 1319 958
rect 1589 543 1800 567
rect 1589 371 1640 543
rect 1752 371 1800 543
rect 1589 346 1800 371
rect 1983 543 2194 572
rect 1983 371 2040 543
rect 2152 371 2194 543
rect 1983 351 2194 371
rect 748 230 819 248
rect 748 197 762 230
rect 804 197 819 230
rect 748 180 819 197
rect 892 180 941 248
rect 679 117 707 118
rect 272 83 707 117
rect 678 82 707 83
rect 683 -268 707 82
rect 678 -269 707 -268
rect 893 -269 941 180
rect 678 -276 711 -269
rect 860 -290 941 -269
rect 989 -341 1028 313
rect 1159 308 1335 333
rect 1159 177 1193 308
rect 1306 177 1335 308
rect 1159 152 1335 177
rect -159 -410 33 -368
rect 817 -409 1028 -341
rect -885 -555 -702 -522
rect -441 -614 -265 -589
rect -441 -745 -407 -614
rect -294 -745 -265 -614
rect 148 -621 295 -509
rect 558 -621 708 -507
rect -441 -771 -265 -745
<< via1 >>
rect 1640 2607 1752 2727
rect 2040 2607 2152 2727
rect -1256 2146 -1131 2319
rect -856 2146 -731 2319
rect 412 2014 480 2076
rect 433 1811 485 1851
rect 1640 1728 1752 1848
rect 2040 1728 2152 1848
rect -1256 1240 -1131 1413
rect -856 1240 -731 1413
rect -375 1009 -315 1018
rect -375 964 -368 1009
rect -368 964 -322 1009
rect -322 964 -315 1009
rect -375 958 -315 964
rect -407 147 -294 266
rect -1256 -522 -1131 -349
rect -856 -522 -731 -349
rect 193 964 221 991
rect 619 1005 650 1007
rect 619 980 620 1005
rect 620 980 648 1005
rect 648 980 650 1005
rect 619 978 650 980
rect 145 770 180 773
rect 145 741 147 770
rect 147 741 178 770
rect 178 741 180 770
rect 145 739 180 741
rect 650 739 695 776
rect 48 227 90 230
rect 48 200 51 227
rect 51 200 87 227
rect 87 200 90 227
rect 48 197 90 200
rect 1640 1122 1752 1242
rect 2040 1122 2152 1242
rect 1225 1009 1285 1018
rect 1225 964 1232 1009
rect 1232 964 1278 1009
rect 1278 964 1285 1009
rect 1225 958 1285 964
rect 1640 371 1752 543
rect 2040 371 2152 543
rect 762 227 804 230
rect 762 200 765 227
rect 765 200 801 227
rect 801 200 804 227
rect 762 197 804 200
rect 1193 192 1306 308
rect 1193 177 1305 192
rect -407 -745 -294 -614
rect 406 -558 455 -514
<< metal2 >>
rect 1590 2727 2192 2778
rect 1590 2607 1640 2727
rect 1752 2607 2040 2727
rect 2152 2607 2192 2727
rect 1590 2505 2192 2607
rect -1285 2319 -1102 2342
rect -1285 2146 -1256 2319
rect -1131 2146 -1102 2319
rect -1285 2113 -1102 2146
rect -885 2319 -702 2342
rect -885 2146 -856 2319
rect -731 2146 -702 2319
rect -885 2113 -702 2146
rect 381 2086 509 2111
rect 381 2003 401 2086
rect 490 2003 509 2086
rect 381 1984 509 2003
rect 402 1851 516 1859
rect 402 1811 433 1851
rect 485 1843 516 1851
rect 1587 1848 2192 2505
rect 1587 1843 1640 1848
rect 485 1811 1640 1843
rect 402 1810 1640 1811
rect 402 1801 516 1810
rect 1587 1728 1640 1810
rect 1752 1728 2040 1848
rect 2152 1728 2192 1848
rect -1285 1413 -1102 1438
rect -1285 1240 -1256 1413
rect -1131 1240 -1102 1413
rect -1285 1207 -1102 1240
rect -885 1413 -702 1438
rect -885 1240 -856 1413
rect -731 1240 -702 1413
rect -885 1207 -702 1240
rect 1587 1242 2192 1728
rect 1587 1122 1640 1242
rect 1752 1122 2040 1242
rect 2152 1122 2192 1242
rect -419 1036 -281 1056
rect -419 941 -395 1036
rect -299 1011 -281 1036
rect 1181 1036 1319 1056
rect 1181 1022 1205 1036
rect 886 1019 1205 1022
rect 615 1016 1205 1019
rect -299 1000 -251 1011
rect 610 1007 1205 1016
rect -299 991 226 1000
rect -299 964 193 991
rect 221 964 226 991
rect 610 978 619 1007
rect 650 978 1205 1007
rect 610 977 1107 978
rect 610 973 655 977
rect -299 959 226 964
rect -299 958 193 959
rect -299 941 -281 958
rect -419 919 -281 941
rect 1181 941 1205 978
rect 1301 941 1319 1036
rect 1181 919 1319 941
rect 133 773 194 783
rect 133 739 145 773
rect 180 739 194 773
rect 133 729 194 739
rect 641 776 702 790
rect 641 739 650 776
rect 695 739 702 776
rect 641 736 702 739
rect -463 625 -254 702
rect -463 591 -253 625
rect 148 591 178 729
rect -463 542 178 591
rect 658 588 690 736
rect 1587 716 2192 1122
rect 1137 588 1342 699
rect -463 519 -253 542
rect 658 539 1342 588
rect -463 266 -254 519
rect 1137 309 1342 539
rect 1587 543 2194 716
rect 1587 371 1640 543
rect 1752 371 2040 543
rect 2152 371 2194 543
rect -463 147 -407 266
rect -294 240 -254 266
rect 1139 308 1340 309
rect 34 240 104 248
rect -294 230 104 240
rect -294 197 48 230
rect 90 197 104 230
rect -294 187 104 197
rect -294 147 -254 187
rect 34 180 104 187
rect 748 241 818 248
rect 1139 241 1193 308
rect 748 230 1193 241
rect 748 197 762 230
rect 804 197 1193 230
rect 748 187 1193 197
rect 1306 192 1340 308
rect 748 180 818 187
rect -463 42 -254 147
rect 1139 177 1193 187
rect 1305 177 1340 192
rect 1587 180 2194 371
rect -1285 -349 -1102 -324
rect -1285 -522 -1256 -349
rect -1131 -522 -1102 -349
rect -1285 -555 -1102 -522
rect -885 -349 -702 -324
rect -885 -522 -856 -349
rect -731 -522 -702 -349
rect -885 -555 -702 -522
rect -460 -586 -259 42
rect 1139 1 1340 177
rect 1589 83 2194 180
rect 1138 -281 1341 1
rect 397 -514 464 -508
rect 397 -558 406 -514
rect 455 -558 464 -514
rect -460 -614 -258 -586
rect -460 -745 -407 -614
rect -294 -668 -258 -614
rect 397 -668 464 -558
rect -294 -713 465 -668
rect -294 -745 -258 -713
rect 1139 -744 1340 -281
rect -460 -770 -258 -745
rect -460 -831 -259 -770
rect 1140 -831 1340 -744
rect 1590 -629 2192 83
rect -460 -842 -258 -831
rect -460 -843 -256 -842
rect 1140 -843 1341 -831
rect -460 -965 1341 -843
rect 1590 -965 2193 -629
<< via2 >>
rect 1640 2607 1752 2727
rect 2040 2607 2152 2727
rect -1256 2146 -1131 2319
rect -856 2146 -731 2319
rect 401 2076 490 2086
rect 401 2014 412 2076
rect 412 2014 480 2076
rect 480 2014 490 2076
rect 401 2003 490 2014
rect 1640 1728 1752 1848
rect 2040 1728 2152 1848
rect -1256 1240 -1131 1413
rect -856 1240 -731 1413
rect 1640 1122 1752 1242
rect 2040 1122 2152 1242
rect -395 1018 -299 1036
rect -395 958 -375 1018
rect -375 958 -315 1018
rect -315 958 -299 1018
rect 1205 1018 1301 1036
rect -395 941 -299 958
rect 1205 958 1225 1018
rect 1225 958 1285 1018
rect 1285 958 1301 1018
rect 1205 941 1301 958
rect 1640 371 1752 543
rect 2040 371 2152 543
rect -407 147 -294 266
rect 1193 192 1306 308
rect 1193 177 1305 192
rect -1256 -522 -1131 -349
rect -856 -522 -731 -349
rect -407 -745 -294 -614
<< metal3 >>
rect 1605 2727 1783 2757
rect 1605 2607 1640 2727
rect 1752 2607 1783 2727
rect 1605 2574 1783 2607
rect 2004 2727 2183 2757
rect 2004 2607 2040 2727
rect 2152 2607 2183 2727
rect 2004 2574 2183 2607
rect -1285 2319 -1102 2342
rect -1285 2146 -1256 2319
rect -1131 2146 -1102 2319
rect -1285 2113 -1102 2146
rect -885 2319 -702 2342
rect -885 2146 -856 2319
rect -731 2146 -702 2319
rect -885 2113 -702 2146
rect -462 2148 1342 2152
rect -462 2086 1349 2148
rect -462 2003 401 2086
rect 490 2003 1349 2086
rect -462 1971 1349 2003
rect -1285 1413 -1102 1438
rect -1285 1240 -1256 1413
rect -1131 1240 -1102 1413
rect -1285 1207 -1102 1240
rect -885 1413 -702 1438
rect -885 1240 -856 1413
rect -731 1240 -702 1413
rect -885 1207 -702 1240
rect -462 1036 -251 1971
rect -462 941 -395 1036
rect -299 941 -251 1036
rect -462 900 -251 941
rect 1138 1036 1349 1971
rect 1604 1848 1783 1878
rect 1604 1728 1640 1848
rect 1752 1728 1783 1848
rect 1604 1695 1783 1728
rect 2004 1848 2183 1878
rect 2004 1728 2040 1848
rect 2152 1728 2183 1848
rect 2004 1695 2183 1728
rect 1604 1242 1783 1272
rect 1604 1122 1640 1242
rect 1752 1122 1783 1242
rect 1604 1091 1783 1122
rect 2004 1242 2183 1272
rect 2004 1122 2040 1242
rect 2152 1122 2183 1242
rect 2004 1091 2183 1122
rect 1138 941 1205 1036
rect 1301 941 1349 1036
rect 1138 900 1349 941
rect 133 729 194 783
rect 148 727 178 729
rect -461 266 -256 351
rect 1137 309 1342 699
rect 1589 543 1800 567
rect 1589 371 1640 543
rect 1752 371 1800 543
rect 1589 346 1800 371
rect 1983 543 2194 572
rect 1983 371 2040 543
rect 2152 371 2194 543
rect 1983 351 2194 371
rect -461 147 -407 266
rect -294 147 -256 266
rect -461 105 -256 147
rect 1138 308 1342 309
rect 1138 177 1193 308
rect 1306 192 1342 308
rect 1305 177 1342 192
rect -456 101 -259 105
rect 1138 -46 1342 177
rect 1138 -246 1341 -46
rect -1285 -349 -1102 -324
rect -1285 -522 -1256 -349
rect -1131 -522 -1102 -349
rect -1285 -555 -1102 -522
rect -885 -349 -702 -324
rect -885 -522 -856 -349
rect -731 -522 -702 -349
rect -885 -555 -702 -522
rect -461 -614 -258 -520
rect -462 -745 -407 -614
rect -294 -745 -258 -614
rect 1138 -618 1342 -246
rect 1138 -741 1341 -618
rect 1138 -744 1342 -741
rect -462 -842 -258 -745
rect -462 -843 -256 -842
rect 1140 -843 1342 -744
rect -462 -886 1342 -843
rect -460 -965 1342 -886
<< via3 >>
rect 1640 2607 1752 2727
rect 2040 2607 2152 2727
rect -1256 2146 -1131 2319
rect -856 2146 -731 2319
rect -1256 1240 -1131 1413
rect -856 1240 -731 1413
rect 1640 1728 1752 1848
rect 2040 1728 2152 1848
rect 1640 1122 1752 1242
rect 2040 1122 2152 1242
rect 1640 371 1752 543
rect 2040 371 2152 543
rect -1256 -522 -1131 -349
rect -856 -522 -731 -349
<< metal4 >>
rect 1588 2727 2195 2778
rect 1588 2675 1640 2727
rect 1590 2607 1640 2675
rect 1752 2607 2040 2727
rect 2152 2607 2195 2727
rect 1590 2527 2195 2607
rect 1589 2505 2195 2527
rect 1587 2389 2195 2505
rect -1285 2319 -1102 2342
rect -1285 2146 -1256 2319
rect -1131 2146 -1102 2319
rect -1285 2113 -1102 2146
rect -885 2319 -702 2342
rect -885 2146 -856 2319
rect -731 2146 -702 2319
rect -885 2113 -702 2146
rect 1587 1848 2192 2389
rect 1587 1728 1640 1848
rect 1752 1728 2040 1848
rect 2152 1728 2192 1848
rect -1285 1413 -1102 1438
rect -1285 1240 -1256 1413
rect -1131 1240 -1102 1413
rect -1285 1207 -1102 1240
rect -885 1413 -702 1438
rect -885 1240 -856 1413
rect -731 1240 -702 1413
rect -885 1207 -702 1240
rect 1587 1242 2192 1728
rect 1587 1122 1640 1242
rect 1752 1122 2040 1242
rect 2152 1122 2192 1242
rect 1587 716 2192 1122
rect 1587 543 2194 716
rect 1587 371 1640 543
rect 1752 371 2040 543
rect 2152 371 2194 543
rect 1587 180 2194 371
rect 1589 83 2194 180
rect -1285 -349 -1102 -324
rect -1285 -522 -1256 -349
rect -1131 -522 -1102 -349
rect -1285 -555 -1102 -522
rect -885 -349 -702 -324
rect -885 -522 -856 -349
rect -731 -522 -702 -349
rect -885 -555 -702 -522
rect 1590 -629 2192 83
rect 1590 -965 2193 -629
<< via4 >>
rect -1256 2146 -1131 2319
rect -856 2146 -731 2319
rect -1256 1240 -1131 1413
rect -856 1240 -731 1413
rect -1256 -522 -1131 -349
rect -856 -522 -731 -349
<< metal5 >>
rect -1299 2536 -675 2766
rect -1296 2319 -677 2536
rect -1296 2146 -1256 2319
rect -1131 2146 -856 2319
rect -731 2146 -677 2319
rect -1296 1413 -677 2146
rect -1296 1240 -1256 1413
rect -1131 1240 -856 1413
rect -731 1240 -677 1413
rect -1296 1017 -677 1240
rect -1296 535 -673 1017
rect -1296 -349 -677 535
rect -1296 -522 -1256 -349
rect -1131 -522 -856 -349
rect -731 -522 -677 -349
rect -1296 -669 -677 -522
rect -1296 -967 -675 -669
use SR_latch  SR_latch_0 ~/mycomparator_copy1/layout/latch
timestamp 1654337383
transform 1 0 197 0 1 2227
box 0 0 436 474
use latch_3  latch_3_0
timestamp 1654337383
transform 1 0 44 0 1 1319
box -8 0 813 511
use preamp_part12  preamp_part12_0 ~/Documents/Comparator_MPW6/mag/preamp
timestamp 1654337383
transform 1 0 356 0 1 -232
box -360 -330 510 693
use preamp_part22  preamp_part22_0 ~/Documents/Comparator_MPW6/mag/preamp
timestamp 1654337383
transform 1 0 68 0 1 660
box 39 151 658 544
<< labels >>
rlabel poly 483 1945 483 1945 1 CLKBAR
rlabel locali 595 2448 595 2448 3 Outn
rlabel locali 257 2431 257 2431 7 Outp
rlabel metal1 640 -621 640 -621 5 Vp
rlabel metal1 220 -621 220 -621 5 Vn
rlabel metal1 -29 669 -29 669 7 fn
rlabel metal5 -910 -967 -910 -967 5 GND
rlabel metal4 1885 -965 1885 -965 5 VDD
rlabel metal3 395 -965 395 -965 5 CLK
rlabel metal1 1029 2281 1029 2281 3 Dn
rlabel metal1 941 672 941 672 3 fp
rlabel metal1 -159 2279 -159 2279 7 Dp
<< end >>
