magic
tech sky130A
magscale 1 2
timestamp 1651643300
<< nwell >>
rect -720 994 1018 1328
<< poly >>
rect -482 1512 -414 1528
rect -482 1470 -466 1512
rect -430 1470 -414 1512
rect -482 1452 -414 1470
rect 688 1512 756 1528
rect 688 1470 704 1512
rect 744 1470 756 1512
rect 688 1452 756 1470
rect -462 1266 -432 1452
rect 706 1276 738 1452
rect -170 888 -42 908
rect -170 842 -148 888
rect -72 842 -42 888
rect -170 802 -42 842
rect 318 800 348 812
rect 414 798 444 810
rect -168 434 -138 464
rect -72 436 -42 466
rect 220 384 446 462
rect -656 326 -594 342
rect 220 340 298 384
rect -656 284 -640 326
rect -606 284 -594 326
rect -656 268 -594 284
rect 218 336 300 340
rect 218 294 236 336
rect 284 294 300 336
rect -640 242 -610 268
rect 218 266 300 294
rect 864 328 926 344
rect 864 286 880 328
rect 914 286 926 328
rect 864 270 926 286
rect 882 234 912 270
rect -434 4 -404 6
rect -338 4 -308 6
rect -242 4 -212 6
rect -146 4 -116 6
rect -434 -168 -116 4
rect -434 -234 -406 -168
rect -144 -234 -116 -168
rect -434 -260 -116 -234
rect 80 -170 206 58
rect 80 -238 104 -170
rect 180 -238 206 -170
rect 80 -258 206 -238
rect 388 -2 418 4
rect 484 -2 514 4
rect 580 -2 610 4
rect 676 -2 706 4
rect 388 -164 706 -2
rect 388 -234 414 -164
rect 680 -234 706 -164
rect 388 -260 706 -234
<< polycont >>
rect -466 1470 -430 1512
rect 704 1470 744 1512
rect -148 842 -72 888
rect -640 284 -606 326
rect 236 294 284 336
rect 880 286 914 328
rect -406 -234 -144 -168
rect 104 -238 180 -170
rect 414 -234 680 -164
<< locali >>
rect -482 1512 -414 1528
rect -482 1470 -466 1512
rect -430 1470 -414 1512
rect -482 1452 -414 1470
rect 688 1512 756 1528
rect 688 1470 704 1512
rect 744 1470 756 1512
rect 688 1452 756 1470
rect -720 1336 1020 1386
rect -508 1208 -474 1336
rect 748 1210 782 1336
rect -164 896 -56 904
rect -164 832 -158 896
rect -60 832 -56 896
rect -164 826 -56 832
rect -218 434 -184 748
rect -26 434 8 746
rect 268 434 302 742
rect 460 434 494 739
rect -218 392 100 434
rect 180 392 494 434
rect -656 326 -594 342
rect -656 284 -642 326
rect -606 284 -594 326
rect -418 312 -412 350
rect -352 340 298 352
rect -352 336 300 340
rect -352 312 236 336
rect -418 308 236 312
rect -418 306 -352 308
rect -656 268 -594 284
rect 218 294 236 308
rect 284 294 300 336
rect -484 238 -66 272
rect 218 266 300 294
rect 864 328 926 344
rect 864 286 878 328
rect 914 286 926 328
rect -718 44 -652 200
rect -484 188 -450 238
rect -292 194 -258 238
rect -100 190 -66 238
rect 338 238 756 272
rect 864 270 926 286
rect 338 192 372 238
rect 530 194 564 238
rect 722 192 756 238
rect -598 -22 -564 52
rect 30 48 66 88
rect 122 87 166 148
rect 222 48 256 86
rect 30 -22 256 48
rect 836 -22 870 54
rect 954 42 1020 198
rect -720 -74 1020 -22
rect -422 -166 -128 -150
rect -422 -234 -406 -166
rect -144 -234 -128 -166
rect -422 -252 -128 -234
rect 78 -170 206 -152
rect 78 -238 104 -170
rect 180 -238 206 -170
rect 78 -260 206 -238
rect 398 -164 696 -148
rect 398 -234 414 -164
rect 680 -234 696 -164
rect 398 -250 696 -234
<< viali >>
rect -466 1470 -430 1512
rect 704 1470 744 1512
rect -158 888 -60 896
rect -158 842 -148 888
rect -148 842 -72 888
rect -72 842 -60 888
rect -158 832 -60 842
rect 100 386 180 434
rect -642 284 -640 326
rect -640 284 -606 326
rect -412 312 -352 350
rect 878 286 880 328
rect 880 286 914 328
rect -406 -168 -144 -166
rect -406 -234 -144 -168
rect 106 -238 180 -170
rect 414 -234 680 -164
<< metal1 >>
rect -482 1512 -414 1528
rect -482 1470 -466 1512
rect -430 1470 -414 1512
rect -482 1452 -414 1470
rect 688 1512 756 1528
rect 688 1470 704 1512
rect 744 1470 756 1512
rect 688 1452 756 1470
rect -428 362 -380 1104
rect -170 896 -46 910
rect -170 832 -158 896
rect -60 886 -46 896
rect 654 886 702 1132
rect -60 838 702 886
rect -60 832 -46 838
rect -170 818 -46 832
rect -428 350 -346 362
rect -656 326 -594 342
rect -428 326 -412 350
rect -718 284 -642 326
rect -606 312 -412 326
rect -352 330 -346 350
rect -352 312 -160 330
rect -606 284 -160 312
rect -656 268 -594 284
rect -692 190 -648 212
rect -390 154 -352 284
rect -198 150 -160 284
rect -122 272 -88 668
rect 88 434 194 450
rect 88 386 100 434
rect 180 386 194 434
rect 88 372 194 386
rect -128 236 -66 272
rect -104 138 -66 236
rect 120 116 166 372
rect 364 272 398 536
rect 654 326 702 838
rect 864 328 926 344
rect 864 326 878 328
rect 434 286 878 326
rect 914 326 926 328
rect 914 286 1020 326
rect 434 284 1020 286
rect 338 238 406 272
rect 338 180 374 238
rect 434 188 470 284
rect 624 192 660 284
rect 864 270 926 284
rect -422 -166 -128 -150
rect -422 -234 -406 -166
rect -144 -234 -128 -166
rect -422 -254 -128 -234
rect 78 -170 206 -152
rect 78 -238 106 -170
rect 180 -238 206 -170
rect 78 -258 206 -238
rect 398 -164 696 -148
rect 398 -234 414 -164
rect 680 -234 696 -164
rect 398 -250 696 -234
use sky130_fd_pr__nfet_01v8_8FHE5N  sky130_fd_pr__nfet_01v8_8FHE5N_0
timestamp 1646423143
transform 1 0 143 0 1 126
box -125 -76 125 76
use sky130_fd_pr__nfet_01v8_F5U58G#1  sky130_fd_pr__nfet_01v8_F5U58G_0
timestamp 1646431323
transform 1 0 -625 0 1 116
box -73 -126 73 126
use sky130_fd_pr__nfet_01v8_F5U58G#1  sky130_fd_pr__nfet_01v8_F5U58G_1
timestamp 1646431323
transform 1 0 897 0 1 120
box -73 -126 73 126
use sky130_fd_pr__nfet_01v8_G6PLX8  sky130_fd_pr__nfet_01v8_G6PLX8_0
timestamp 1646422066
transform 1 0 -275 0 1 122
box -221 -126 221 150
use sky130_fd_pr__nfet_01v8_G6PLX8  sky130_fd_pr__nfet_01v8_G6PLX8_1
timestamp 1646422066
transform 1 0 547 0 1 122
box -221 -126 221 150
use sky130_fd_pr__nfet_01v8_RURP52  sky130_fd_pr__nfet_01v8_RURP52_0
timestamp 1651643300
transform 1 0 -105 0 1 630
box -125 -176 125 176
use sky130_fd_pr__nfet_01v8_RURP52  sky130_fd_pr__nfet_01v8_RURP52_1
timestamp 1651643300
transform 1 0 381 0 1 630
box -125 -176 125 176
use sky130_fd_pr__pfet_01v8_RFM3CD#0  sky130_fd_pr__pfet_01v8_RFM3CD_0
timestamp 1646431323
transform 1 0 -447 0 1 1160
box -109 -162 109 162
use sky130_fd_pr__pfet_01v8_RFM3CD#0  sky130_fd_pr__pfet_01v8_RFM3CD_1
timestamp 1646431323
transform 1 0 721 0 1 1160
box -109 -162 109 162
<< end >>
