* SPICE3 file created from user_analog_project_wrapper.ext - technology: sky130A

.subckt sky130_fd_pr__diode_pw2nd_05v5_3P6M5Y a_n100_n100# w_n238_n238#
D0 w_n238_n238# a_n100_n100# sky130_fd_pr__diode_pw2nd_05v5 pj=4e+06u area=1e+12p
.ends

.subckt sky130_fd_pr__diode_pd2nw_05v5_RT56W3 w_n321_n321# a_n45_n45# w_n183_n183#
D0 a_n45_n45# w_n183_n183# sky130_fd_pr__diode_pd2nw_05v5 pj=1.8e+06u area=2.025e+11p
.ends

.subckt sky130_fd_sc_hd__buf_2 A VGND VPWR X VNB VPB
X0 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=5.63e+11p pd=5.18e+06u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X1 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X3 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=3.6625e+11p ps=3.78e+06u w=650000u l=150000u
X4 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
.ends

.subckt sky130_fd_sc_hd__buf_16 A VGND VPWR X VNB VPB
X0 VGND A a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=2.093e+12p pd=2.204e+07u as=5.265e+11p ps=5.52e+06u w=650000u l=150000u
X1 X a_109_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=2.16e+12p pd=2.032e+07u as=3.22e+12p ps=3.044e+07u w=1e+06u l=150000u
X2 VGND a_109_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.404e+12p ps=1.472e+07u w=650000u l=150000u
X3 VGND a_109_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 X a_109_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 VGND a_109_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 VPWR a_109_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 a_109_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=8.1e+11p pd=7.62e+06u as=0p ps=0u w=1e+06u l=150000u
X8 X a_109_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 VPWR A a_109_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 X a_109_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 X a_109_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 X a_109_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 X a_109_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X14 a_109_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 VPWR a_109_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16 X a_109_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X17 X a_109_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X18 VPWR A a_109_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X19 VPWR a_109_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X20 VGND A a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X21 VGND A a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X22 VGND a_109_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X23 X a_109_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X24 VGND a_109_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X25 VPWR a_109_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X26 VGND a_109_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X27 VPWR a_109_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X28 X a_109_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X29 VGND a_109_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X30 a_109_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X31 a_109_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X32 X a_109_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X33 VPWR a_109_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X34 X a_109_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X35 X a_109_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X36 VPWR A a_109_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X37 X a_109_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X38 X a_109_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X39 a_109_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X40 VPWR a_109_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X41 VPWR a_109_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X42 a_109_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X43 VGND a_109_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
C0 X VPWR 3.72fF
C1 X VGND 2.53fF
C2 X a_109_47# 4.49fF
C3 VPWR VPB 2.24fF
C4 VPB VNB 2.02fF
.ends

.subckt sky130_fd_pr__diode_pw2nd_05v5_GT7G3L a_n45_n45# w_n183_n183#
D0 w_n183_n183# a_n45_n45# sky130_fd_pr__diode_pw2nd_05v5 pj=1.8e+06u area=2.025e+11p
.ends

.subckt sky130_fd_pr__pfet_01v8_GJYUB2 a_207_n100# a_81_n126# a_n207_n128# a_15_n100#
+ a_n177_n100# a_111_n100# a_n15_n128# a_n111_n126# w_n305_n200# a_n81_n100# a_177_n128#
+ a_n269_n100# VSUBS
X0 a_207_n100# a_177_n128# a_111_n100# w_n305_n200# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.3e+11p ps=2.66e+06u w=1e+06u l=150000u
X1 a_15_n100# a_n15_n128# a_n81_n100# w_n305_n200# sky130_fd_pr__pfet_01v8 ad=3.3e+11p pd=2.66e+06u as=3.3e+11p ps=2.66e+06u w=1e+06u l=150000u
X2 a_111_n100# a_81_n126# a_15_n100# w_n305_n200# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 a_n81_n100# a_n111_n126# a_n177_n100# w_n305_n200# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=3.3e+11p ps=2.66e+06u w=1e+06u l=150000u
X4 a_n177_n100# a_n207_n128# a_n269_n100# w_n305_n200# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
.ends

.subckt sky130_fd_pr__nfet_01v8_7RYEVP a_n73_n69# a_n15_n89# a_15_n69# VSUBS
X0 a_15_n69# a_n15_n89# a_n73_n69# VSUBS sky130_fd_pr__nfet_01v8 ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=150000u
.ends

.subckt nmos_1u#0 sky130_fd_pr__nfet_01v8_7RYEVP_0/a_n15_n89# sky130_fd_pr__nfet_01v8_7RYEVP_0/a_15_n69#
+ sky130_fd_pr__nfet_01v8_7RYEVP_0/a_n73_n69# VSUBS
Xsky130_fd_pr__nfet_01v8_7RYEVP_0 sky130_fd_pr__nfet_01v8_7RYEVP_0/a_n73_n69# sky130_fd_pr__nfet_01v8_7RYEVP_0/a_n15_n89#
+ sky130_fd_pr__nfet_01v8_7RYEVP_0/a_15_n69# VSUBS sky130_fd_pr__nfet_01v8_7RYEVP
.ends

.subckt pmos_2uf2#0 a_n139_n100# a_63_n100# a_33_n130# a_n33_n100# w_n319_n202# a_n63_n130#
+ VSUBS
X0 a_63_n100# a_33_n130# a_n33_n100# w_n319_n202# sky130_fd_pr__pfet_01v8 ad=3.048e+11p pd=2.62e+06u as=3.3e+11p ps=2.66e+06u w=1e+06u l=150000u
X1 a_n33_n100# a_n63_n130# a_n139_n100# w_n319_n202# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=3.8e+11p ps=2.76e+06u w=1e+06u l=150000u
.ends

.subckt inv_W12 Vout Vin VDD GND pmos_2uf2_0/w_n319_n202# nmos_1u_0/sky130_fd_pr__nfet_01v8_7RYEVP_0/a_15_n69#
+ VSUBS
Xnmos_1u_0 Vin nmos_1u_0/sky130_fd_pr__nfet_01v8_7RYEVP_0/a_15_n69# GND VSUBS nmos_1u#0
Xpmos_2uf2_0 VDD VDD Vin Vout pmos_2uf2_0/w_n319_n202# Vin VSUBS pmos_2uf2#0
.ends

.subckt latch_3 a_646_808# inv_W12_1/GND m1_686_734# w_n16_492# inv_W12_1/Vin VSUBS
+ inv_W12_0/Vin
Xsky130_fd_pr__pfet_01v8_GJYUB2_0 m1_686_734# a_646_808# a_646_808# m1_686_734# m1_686_734#
+ inv_W12_1/VDD a_646_808# a_646_808# w_n16_492# inv_W12_1/VDD a_646_808# inv_W12_1/VDD
+ VSUBS sky130_fd_pr__pfet_01v8_GJYUB2
Xinv_W12_0 inv_W12_1/Vin inv_W12_0/Vin inv_W12_1/VDD inv_W12_1/GND w_n16_492# inv_W12_1/Vin
+ VSUBS inv_W12
Xinv_W12_1 inv_W12_0/Vin inv_W12_1/Vin inv_W12_1/VDD inv_W12_1/GND w_n16_492# inv_W12_0/Vin
+ VSUBS inv_W12
C0 w_n16_492# VSUBS 2.44fF
.ends

.subckt sky130_fd_pr__nfet_01v8_G6PLX8 a_n129_n500# a_63_n500# a_n221_n474# a_n33_n500#
+ a_n159_n522# a_159_n500# VSUBS
X0 a_n33_n500# a_n159_n522# a_n129_n500# VSUBS sky130_fd_pr__nfet_01v8 ad=3.3e+11p pd=2.66e+06u as=3.3e+11p ps=2.66e+06u w=1e+06u l=150000u
X1 a_159_n500# a_n159_n522# a_63_n500# VSUBS sky130_fd_pr__nfet_01v8 ad=3.048e+11p pd=2.62e+06u as=3.3e+11p ps=2.66e+06u w=1e+06u l=150000u
X2 a_63_n500# a_n159_n522# a_n33_n500# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 a_n129_n500# a_n159_n522# a_n221_n474# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.048e+11p ps=2.62e+06u w=1e+06u l=150000u
.ends

.subckt sky130_fd_pr__pfet_01v8_RFM3CD#0 a_n73_n100# w_n109_n162# a_15_n100# a_n15_n126#
+ VSUBS
X0 a_15_n100# a_n15_n126# a_n73_n100# w_n109_n162# sky130_fd_pr__pfet_01v8 ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=150000u
.ends

.subckt sky130_fd_pr__nfet_01v8_F5U58G#1 a_15_n500# a_n15_n526# a_n73_n500# VSUBS
X0 a_15_n500# a_n15_n526# a_n73_n500# VSUBS sky130_fd_pr__nfet_01v8 ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=150000u
.ends

.subckt sky130_fd_pr__nfet_01v8_RURP52 a_33_n370# a_63_n348# a_n63_n370# a_n33_n348#
+ a_n125_n348# VSUBS
X0 a_n33_n348# a_n63_n370# a_n125_n348# VSUBS sky130_fd_pr__nfet_01v8 ad=4.95e+11p pd=3.66e+06u as=4.65e+11p ps=3.62e+06u w=1.5e+06u l=150000u
X1 a_63_n348# a_33_n370# a_n33_n348# VSUBS sky130_fd_pr__nfet_01v8 ad=4.65e+11p pd=3.62e+06u as=0p ps=0u w=1.5e+06u l=150000u
.ends

.subckt sky130_fd_pr__nfet_01v8_8FHE5N a_n125_n439# a_63_n450# a_n63_n476# a_n33_n450#
+ a_33_n476# VSUBS
X0 a_63_n450# a_33_n476# a_n33_n450# VSUBS sky130_fd_pr__nfet_01v8 ad=1.528e+11p pd=1.62e+06u as=1.65e+11p ps=1.66e+06u w=500000u l=150000u
X1 a_n33_n450# a_n63_n476# a_n125_n439# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.528e+11p ps=1.62e+06u w=500000u l=150000u
.ends

.subckt preamp_part12 li_n720_1336# a_n72_236# a_80_n658# a_n434_n660# m1_n692_n210#
+ a_n506_870# a_388_n660# w_n720_994# li_n720_n474# a_414_256# a_706_862# li_954_n358#
+ VSUBS
Xsky130_fd_pr__nfet_01v8_G6PLX8_0 a_414_256# a_414_256# m1_n128_n164# m1_n128_n164#
+ a_n434_n660# m1_n128_n164# VSUBS sky130_fd_pr__nfet_01v8_G6PLX8
Xsky130_fd_pr__nfet_01v8_G6PLX8_1 a_n72_236# a_n72_236# m1_338_n220# m1_338_n220#
+ a_388_n660# m1_338_n220# VSUBS sky130_fd_pr__nfet_01v8_G6PLX8
Xsky130_fd_pr__pfet_01v8_RFM3CD_0 li_n720_1336# w_n720_994# a_414_256# a_n506_870#
+ VSUBS sky130_fd_pr__pfet_01v8_RFM3CD#0
Xsky130_fd_pr__pfet_01v8_RFM3CD_1 a_n72_236# w_n720_994# li_n720_1336# a_706_862#
+ VSUBS sky130_fd_pr__pfet_01v8_RFM3CD#0
Xsky130_fd_pr__nfet_01v8_F5U58G_0 li_n720_n474# a_414_256# m1_n692_n210# VSUBS sky130_fd_pr__nfet_01v8_F5U58G#1
Xsky130_fd_pr__nfet_01v8_F5U58G_1 li_954_n358# a_n72_236# li_n720_n474# VSUBS sky130_fd_pr__nfet_01v8_F5U58G#1
Xsky130_fd_pr__nfet_01v8_RURP52_0 a_n72_236# li_n218_192# a_n72_236# m1_n128_n164#
+ li_n218_192# VSUBS sky130_fd_pr__nfet_01v8_RURP52
Xsky130_fd_pr__nfet_01v8_RURP52_1 a_414_256# li_n218_192# a_414_256# m1_338_n220#
+ li_n218_192# VSUBS sky130_fd_pr__nfet_01v8_RURP52
Xsky130_fd_pr__nfet_01v8_8FHE5N_0 li_n720_n474# li_n720_n474# a_80_n658# li_n218_192#
+ a_80_n658# VSUBS sky130_fd_pr__nfet_01v8_8FHE5N
C0 w_n720_994# VSUBS 2.08fF
.ends

.subckt sky130_fd_pr__nfet_01v8_F5U58G a_n73_n100# a_15_n100# a_n15_n126# VSUBS
X0 a_15_n100# a_n15_n126# a_n73_n100# VSUBS sky130_fd_pr__nfet_01v8 ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=150000u
.ends

.subckt sky130_fd_pr__pfet_01v8_AC5E9B w_n161_n200# a_33_n126# a_63_n100# a_n125_n74#
+ a_n33_n100# a_n63_n130# VSUBS
X0 a_63_n100# a_33_n126# a_n33_n100# w_n161_n200# sky130_fd_pr__pfet_01v8 ad=3.048e+11p pd=2.62e+06u as=3.3e+11p ps=2.66e+06u w=1e+06u l=150000u
X1 a_n33_n100# a_n63_n130# a_n125_n74# w_n161_n200# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=3.048e+11p ps=2.62e+06u w=1e+06u l=150000u
.ends

.subckt SR_latch a_648_848# sky130_fd_pr__nfet_01v8_F5U58G_1/a_n15_n126# sky130_fd_pr__nfet_01v8_F5U58G_0/a_n15_n126#
+ a_262_508# VDD w_0_524# GND VSUBS
Xsky130_fd_pr__nfet_01v8_F5U58G_0 a_648_848# GND sky130_fd_pr__nfet_01v8_F5U58G_0/a_n15_n126#
+ VSUBS sky130_fd_pr__nfet_01v8_F5U58G
Xsky130_fd_pr__nfet_01v8_F5U58G_1 GND a_262_508# sky130_fd_pr__nfet_01v8_F5U58G_1/a_n15_n126#
+ VSUBS sky130_fd_pr__nfet_01v8_F5U58G
Xsky130_fd_pr__pfet_01v8_AC5E9B_0 w_0_524# a_262_508# VDD VDD a_648_848# a_262_508#
+ VSUBS sky130_fd_pr__pfet_01v8_AC5E9B
Xsky130_fd_pr__pfet_01v8_AC5E9B_1 w_0_524# a_648_848# VDD VDD a_262_508# a_648_848#
+ VSUBS sky130_fd_pr__pfet_01v8_AC5E9B
.ends

.subckt preamp_part22 w_78_306# a_392_716# sky130_fd_pr__pfet_01v8_RFM3CD#0_0/a_n15_n126#
+ sky130_fd_pr__pfet_01v8_RFM3CD#0_1/a_n15_n126# sky130_fd_pr__pfet_01v8_RFM3CD#0_2/a_n15_n126#
+ sky130_fd_pr__pfet_01v8_RFM3CD#0_3/a_n15_n126# a_810_594# li_116_1034# sky130_fd_pr__pfet_01v8_RFM3CD#0_3/a_15_n100#
+ VSUBS sky130_fd_pr__pfet_01v8_RFM3CD#0_2/a_n73_n100#
Xsky130_fd_pr__pfet_01v8_RFM3CD#0_0 li_214_402# w_78_306# a_810_594# sky130_fd_pr__pfet_01v8_RFM3CD#0_0/a_n15_n126#
+ VSUBS sky130_fd_pr__pfet_01v8_RFM3CD#0
Xsky130_fd_pr__pfet_01v8_RFM3CD#0_1 a_392_716# w_78_306# li_1016_536# sky130_fd_pr__pfet_01v8_RFM3CD#0_1/a_n15_n126#
+ VSUBS sky130_fd_pr__pfet_01v8_RFM3CD#0
Xsky130_fd_pr__pfet_01v8_RFM3CD#0_2 sky130_fd_pr__pfet_01v8_RFM3CD#0_2/a_n73_n100#
+ w_78_306# li_214_402# sky130_fd_pr__pfet_01v8_RFM3CD#0_2/a_n15_n126# VSUBS sky130_fd_pr__pfet_01v8_RFM3CD#0
Xsky130_fd_pr__pfet_01v8_RFM3CD#0_3 li_1016_536# w_78_306# sky130_fd_pr__pfet_01v8_RFM3CD#0_3/a_15_n100#
+ sky130_fd_pr__pfet_01v8_RFM3CD#0_3/a_n15_n126# VSUBS sky130_fd_pr__pfet_01v8_RFM3CD#0
Xsky130_fd_pr__pfet_01v8_RFM3CD_0 li_214_402# w_78_306# li_116_1034# a_392_716# VSUBS
+ sky130_fd_pr__pfet_01v8_RFM3CD#0
Xsky130_fd_pr__pfet_01v8_RFM3CD_1 li_116_1034# w_78_306# li_1016_536# a_810_594# VSUBS
+ sky130_fd_pr__pfet_01v8_RFM3CD#0
C0 w_78_306# VSUBS 2.70fF
.ends

.subckt comparator_v6 Outn Vp Vn CLK VDD GND Outp CLKBAR
Xlatch_3_0 CLKBAR GND VDD VDD Dp GND Dn latch_3
Xpreamp_part12_0 VDD fp CLK Vn Dp CLK Vp VDD GND fn CLK Dn GND preamp_part12
XSR_latch_0 Outp Dn Dp Outn VDD VDD GND GND SR_latch
Xpreamp_part22_0 VDD fp CLKBAR CLKBAR CLK CLK fn VDD VDD GND VDD preamp_part22
C0 VDD CLKBAR 2.34fF
C1 VDD GND 29.75fF
C2 CLK GND 14.11fF
C3 fp GND 2.32fF
C4 fn GND 2.31fF
C5 Dp GND 3.77fF
C6 Dn GND 3.24fF
C7 CLKBAR GND 3.04fF
.ends

.subckt user_analog_project_wrapper gpio_analog[0] gpio_analog[10] gpio_analog[11]
+ gpio_analog[12] gpio_analog[13] gpio_analog[14] gpio_analog[15] gpio_analog[16]
+ gpio_analog[17] gpio_analog[1] gpio_analog[2] gpio_analog[3] gpio_analog[4] gpio_analog[5]
+ gpio_analog[6] gpio_analog[7] gpio_analog[8] gpio_analog[9] gpio_noesd[0] gpio_noesd[10]
+ gpio_noesd[11] gpio_noesd[12] gpio_noesd[13] gpio_noesd[14] gpio_noesd[15] gpio_noesd[16]
+ gpio_noesd[17] gpio_noesd[1] gpio_noesd[2] gpio_noesd[3] gpio_noesd[4] gpio_noesd[5]
+ gpio_noesd[6] gpio_noesd[7] gpio_noesd[8] gpio_noesd[9] io_analog[0] io_analog[10]
+ io_analog[1] io_analog[2] io_analog[3] io_analog[6] io_analog[7] io_analog[8] io_analog[9]
+ io_analog[4] io_analog[5] io_clamp_high[0] io_clamp_high[1] io_clamp_high[2] io_clamp_low[0]
+ io_clamp_low[1] io_clamp_low[2] io_in[0] io_in[10] io_in[11] io_in[12] io_in[13]
+ io_in[14] io_in[15] io_in[16] io_in[17] io_in[18] io_in[19] io_in[1] io_in[20] io_in[21]
+ io_in[22] io_in[23] io_in[24] io_in[25] io_in[26] io_in[2] io_in[3] io_in[4] io_in[5]
+ io_in[6] io_in[7] io_in[8] io_in[9] io_in_3v3[0] io_in_3v3[10] io_in_3v3[11] io_in_3v3[12]
+ io_in_3v3[13] io_in_3v3[14] io_in_3v3[15] io_in_3v3[16] io_in_3v3[17] io_in_3v3[18]
+ io_in_3v3[19] io_in_3v3[1] io_in_3v3[20] io_in_3v3[21] io_in_3v3[22] io_in_3v3[23]
+ io_in_3v3[24] io_in_3v3[25] io_in_3v3[26] io_in_3v3[2] io_in_3v3[3] io_in_3v3[4]
+ io_in_3v3[5] io_in_3v3[6] io_in_3v3[7] io_in_3v3[8] io_in_3v3[9] io_oeb[0] io_oeb[10]
+ io_oeb[11] io_oeb[12] io_oeb[13] io_oeb[14] io_oeb[15] io_oeb[16] io_oeb[17] io_oeb[18]
+ io_oeb[19] io_oeb[1] io_oeb[20] io_oeb[21] io_oeb[22] io_oeb[23] io_oeb[24] io_oeb[25]
+ io_oeb[26] io_oeb[2] io_oeb[3] io_oeb[4] io_oeb[5] io_oeb[6] io_oeb[7] io_oeb[8]
+ io_oeb[9] io_out[0] io_out[10] io_out[11] io_out[12] io_out[13] io_out[14] io_out[15]
+ io_out[16] io_out[17] io_out[18] io_out[19] io_out[1] io_out[20] io_out[21] io_out[22]
+ io_out[23] io_out[24] io_out[25] io_out[26] io_out[2] io_out[3] io_out[4] io_out[5]
+ io_out[6] io_out[7] io_out[8] io_out[9] la_data_in[0] la_data_in[100] la_data_in[101]
+ la_data_in[102] la_data_in[103] la_data_in[104] la_data_in[105] la_data_in[106]
+ la_data_in[107] la_data_in[108] la_data_in[109] la_data_in[10] la_data_in[110] la_data_in[111]
+ la_data_in[112] la_data_in[113] la_data_in[114] la_data_in[115] la_data_in[116]
+ la_data_in[117] la_data_in[118] la_data_in[119] la_data_in[11] la_data_in[120] la_data_in[121]
+ la_data_in[122] la_data_in[123] la_data_in[124] la_data_in[125] la_data_in[126]
+ la_data_in[127] la_data_in[12] la_data_in[13] la_data_in[14] la_data_in[15] la_data_in[16]
+ la_data_in[17] la_data_in[18] la_data_in[19] la_data_in[1] la_data_in[20] la_data_in[21]
+ la_data_in[22] la_data_in[23] la_data_in[24] la_data_in[25] la_data_in[26] la_data_in[27]
+ la_data_in[28] la_data_in[29] la_data_in[2] la_data_in[30] la_data_in[31] la_data_in[32]
+ la_data_in[33] la_data_in[34] la_data_in[35] la_data_in[36] la_data_in[37] la_data_in[38]
+ la_data_in[39] la_data_in[3] la_data_in[40] la_data_in[41] la_data_in[42] la_data_in[43]
+ la_data_in[44] la_data_in[45] la_data_in[46] la_data_in[47] la_data_in[48] la_data_in[49]
+ la_data_in[4] la_data_in[50] la_data_in[51] la_data_in[52] la_data_in[53] la_data_in[54]
+ la_data_in[55] la_data_in[56] la_data_in[57] la_data_in[58] la_data_in[59] la_data_in[5]
+ la_data_in[60] la_data_in[61] la_data_in[62] la_data_in[63] la_data_in[64] la_data_in[65]
+ la_data_in[66] la_data_in[67] la_data_in[68] la_data_in[69] la_data_in[6] la_data_in[70]
+ la_data_in[71] la_data_in[72] la_data_in[73] la_data_in[74] la_data_in[75] la_data_in[76]
+ la_data_in[77] la_data_in[78] la_data_in[79] la_data_in[7] la_data_in[80] la_data_in[81]
+ la_data_in[82] la_data_in[83] la_data_in[84] la_data_in[85] la_data_in[86] la_data_in[87]
+ la_data_in[88] la_data_in[89] la_data_in[8] la_data_in[90] la_data_in[91] la_data_in[92]
+ la_data_in[93] la_data_in[94] la_data_in[95] la_data_in[96] la_data_in[97] la_data_in[98]
+ la_data_in[99] la_data_in[9] la_data_out[0] la_data_out[100] la_data_out[101] la_data_out[102]
+ la_data_out[103] la_data_out[104] la_data_out[105] la_data_out[106] la_data_out[107]
+ la_data_out[108] la_data_out[109] la_data_out[10] la_data_out[110] la_data_out[111]
+ la_data_out[112] la_data_out[113] la_data_out[114] la_data_out[115] la_data_out[116]
+ la_data_out[117] la_data_out[118] la_data_out[119] la_data_out[11] la_data_out[120]
+ la_data_out[121] la_data_out[122] la_data_out[123] la_data_out[124] la_data_out[125]
+ la_data_out[126] la_data_out[127] la_data_out[12] la_data_out[13] la_data_out[14]
+ la_data_out[15] la_data_out[16] la_data_out[17] la_data_out[18] la_data_out[19]
+ la_data_out[1] la_data_out[20] la_data_out[21] la_data_out[22] la_data_out[23] la_data_out[24]
+ la_data_out[25] la_data_out[26] la_data_out[27] la_data_out[28] la_data_out[29]
+ la_data_out[2] la_data_out[30] la_data_out[31] la_data_out[32] la_data_out[33] la_data_out[34]
+ la_data_out[35] la_data_out[36] la_data_out[37] la_data_out[38] la_data_out[39]
+ la_data_out[3] la_data_out[40] la_data_out[41] la_data_out[42] la_data_out[43] la_data_out[44]
+ la_data_out[45] la_data_out[46] la_data_out[47] la_data_out[48] la_data_out[49]
+ la_data_out[4] la_data_out[50] la_data_out[51] la_data_out[52] la_data_out[53] la_data_out[54]
+ la_data_out[55] la_data_out[56] la_data_out[57] la_data_out[58] la_data_out[59]
+ la_data_out[5] la_data_out[60] la_data_out[61] la_data_out[62] la_data_out[63] la_data_out[64]
+ la_data_out[65] la_data_out[66] la_data_out[67] la_data_out[68] la_data_out[69]
+ la_data_out[6] la_data_out[70] la_data_out[71] la_data_out[72] la_data_out[73] la_data_out[74]
+ la_data_out[75] la_data_out[76] la_data_out[77] la_data_out[78] la_data_out[79]
+ la_data_out[7] la_data_out[80] la_data_out[81] la_data_out[82] la_data_out[83] la_data_out[84]
+ la_data_out[85] la_data_out[86] la_data_out[87] la_data_out[88] la_data_out[89]
+ la_data_out[8] la_data_out[90] la_data_out[91] la_data_out[92] la_data_out[93] la_data_out[94]
+ la_data_out[95] la_data_out[96] la_data_out[97] la_data_out[98] la_data_out[99]
+ la_data_out[9] la_oenb[0] la_oenb[100] la_oenb[101] la_oenb[102] la_oenb[103] la_oenb[104]
+ la_oenb[105] la_oenb[106] la_oenb[107] la_oenb[108] la_oenb[109] la_oenb[10] la_oenb[110]
+ la_oenb[111] la_oenb[112] la_oenb[113] la_oenb[114] la_oenb[115] la_oenb[116] la_oenb[117]
+ la_oenb[118] la_oenb[119] la_oenb[11] la_oenb[120] la_oenb[121] la_oenb[122] la_oenb[123]
+ la_oenb[124] la_oenb[125] la_oenb[126] la_oenb[127] la_oenb[12] la_oenb[13] la_oenb[14]
+ la_oenb[15] la_oenb[16] la_oenb[17] la_oenb[18] la_oenb[19] la_oenb[1] la_oenb[20]
+ la_oenb[21] la_oenb[22] la_oenb[23] la_oenb[24] la_oenb[25] la_oenb[26] la_oenb[27]
+ la_oenb[28] la_oenb[29] la_oenb[2] la_oenb[30] la_oenb[31] la_oenb[32] la_oenb[33]
+ la_oenb[34] la_oenb[35] la_oenb[36] la_oenb[37] la_oenb[38] la_oenb[39] la_oenb[3]
+ la_oenb[40] la_oenb[41] la_oenb[42] la_oenb[43] la_oenb[44] la_oenb[45] la_oenb[46]
+ la_oenb[47] la_oenb[48] la_oenb[49] la_oenb[4] la_oenb[50] la_oenb[51] la_oenb[52]
+ la_oenb[53] la_oenb[54] la_oenb[55] la_oenb[56] la_oenb[57] la_oenb[58] la_oenb[59]
+ la_oenb[5] la_oenb[60] la_oenb[61] la_oenb[62] la_oenb[63] la_oenb[64] la_oenb[65]
+ la_oenb[66] la_oenb[67] la_oenb[68] la_oenb[69] la_oenb[6] la_oenb[70] la_oenb[71]
+ la_oenb[72] la_oenb[73] la_oenb[74] la_oenb[75] la_oenb[76] la_oenb[77] la_oenb[78]
+ la_oenb[79] la_oenb[7] la_oenb[80] la_oenb[81] la_oenb[82] la_oenb[83] la_oenb[84]
+ la_oenb[85] la_oenb[86] la_oenb[87] la_oenb[88] la_oenb[89] la_oenb[8] la_oenb[90]
+ la_oenb[91] la_oenb[92] la_oenb[93] la_oenb[94] la_oenb[95] la_oenb[96] la_oenb[97]
+ la_oenb[98] la_oenb[99] la_oenb[9] user_clock2 user_irq[0] user_irq[1] user_irq[2]
+ vccd1 vccd2 vdda1 vdda2 vssa1 vssa2 vssd1 vssd2 wb_clk_i wb_rst_i wbs_ack_o wbs_adr_i[0]
+ wbs_adr_i[10] wbs_adr_i[11] wbs_adr_i[12] wbs_adr_i[13] wbs_adr_i[14] wbs_adr_i[15]
+ wbs_adr_i[16] wbs_adr_i[17] wbs_adr_i[18] wbs_adr_i[19] wbs_adr_i[1] wbs_adr_i[20]
+ wbs_adr_i[21] wbs_adr_i[22] wbs_adr_i[23] wbs_adr_i[24] wbs_adr_i[25] wbs_adr_i[26]
+ wbs_adr_i[27] wbs_adr_i[28] wbs_adr_i[29] wbs_adr_i[2] wbs_adr_i[30] wbs_adr_i[31]
+ wbs_adr_i[3] wbs_adr_i[4] wbs_adr_i[5] wbs_adr_i[6] wbs_adr_i[7] wbs_adr_i[8] wbs_adr_i[9]
+ wbs_cyc_i wbs_dat_i[0] wbs_dat_i[10] wbs_dat_i[11] wbs_dat_i[12] wbs_dat_i[13] wbs_dat_i[14]
+ wbs_dat_i[15] wbs_dat_i[16] wbs_dat_i[17] wbs_dat_i[18] wbs_dat_i[19] wbs_dat_i[1]
+ wbs_dat_i[20] wbs_dat_i[21] wbs_dat_i[22] wbs_dat_i[23] wbs_dat_i[24] wbs_dat_i[25]
+ wbs_dat_i[26] wbs_dat_i[27] wbs_dat_i[28] wbs_dat_i[29] wbs_dat_i[2] wbs_dat_i[30]
+ wbs_dat_i[31] wbs_dat_i[3] wbs_dat_i[4] wbs_dat_i[5] wbs_dat_i[6] wbs_dat_i[7] wbs_dat_i[8]
+ wbs_dat_i[9] wbs_dat_o[0] wbs_dat_o[10] wbs_dat_o[11] wbs_dat_o[12] wbs_dat_o[13]
+ wbs_dat_o[14] wbs_dat_o[15] wbs_dat_o[16] wbs_dat_o[17] wbs_dat_o[18] wbs_dat_o[19]
+ wbs_dat_o[1] wbs_dat_o[20] wbs_dat_o[21] wbs_dat_o[22] wbs_dat_o[23] wbs_dat_o[24]
+ wbs_dat_o[25] wbs_dat_o[26] wbs_dat_o[27] wbs_dat_o[28] wbs_dat_o[29] wbs_dat_o[2]
+ wbs_dat_o[30] wbs_dat_o[31] wbs_dat_o[3] wbs_dat_o[4] wbs_dat_o[5] wbs_dat_o[6]
+ wbs_dat_o[7] wbs_dat_o[8] wbs_dat_o[9] wbs_sel_i[0] wbs_sel_i[1] wbs_sel_i[2] wbs_sel_i[3]
+ wbs_stb_i wbs_we_i
Xsky130_fd_pr__diode_pw2nd_05v5_3P6M5Y_0 io_analog[7] io_clamp_low[1] sky130_fd_pr__diode_pw2nd_05v5_3P6M5Y
Xsky130_fd_pr__diode_pd2nw_05v5_RT56W3_0 io_clamp_low[1] io_analog[8] io_clamp_high[1]
+ sky130_fd_pr__diode_pd2nw_05v5_RT56W3
Xsky130_fd_pr__diode_pd2nw_05v5_RT56W3_1 io_clamp_low[1] io_analog[7] io_clamp_high[1]
+ sky130_fd_pr__diode_pd2nw_05v5_RT56W3
Xsky130_fd_sc_hd__buf_2_0 comparator_v6_0/Outn io_clamp_low[1] io_clamp_high[1] sky130_fd_sc_hd__buf_2_0/X
+ io_clamp_low[1] io_clamp_high[1] sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_16_0 sky130_fd_sc_hd__buf_2_0/X io_clamp_low[1] io_clamp_high[1]
+ io_analog[3] io_clamp_low[1] io_clamp_high[1] sky130_fd_sc_hd__buf_16
Xsky130_fd_pr__diode_pw2nd_05v5_GT7G3L_0 io_analog[8] io_clamp_low[1] sky130_fd_pr__diode_pw2nd_05v5_GT7G3L
Xsky130_fd_sc_hd__buf_2_1 comparator_v6_0/Outp io_clamp_low[1] io_clamp_high[1] sky130_fd_sc_hd__buf_2_1/X
+ io_clamp_low[1] io_clamp_high[1] sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_16_1 sky130_fd_sc_hd__buf_2_1/X io_clamp_low[1] io_clamp_high[1]
+ io_analog[2] io_clamp_low[1] io_clamp_high[1] sky130_fd_sc_hd__buf_16
Xsky130_fd_sc_hd__buf_2_2 io_analog[8] io_clamp_low[1] io_clamp_high[1] sky130_fd_sc_hd__buf_2_2/X
+ io_clamp_low[1] io_clamp_high[1] sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_16_2 sky130_fd_sc_hd__buf_2_3/X io_clamp_low[1] io_clamp_high[1]
+ comparator_v6_0/CLKBAR io_clamp_low[1] io_clamp_high[1] sky130_fd_sc_hd__buf_16
Xsky130_fd_sc_hd__buf_2_3 io_analog[7] io_clamp_low[1] io_clamp_high[1] sky130_fd_sc_hd__buf_2_3/X
+ io_clamp_low[1] io_clamp_high[1] sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_16_3 sky130_fd_sc_hd__buf_2_2/X io_clamp_low[1] io_clamp_high[1]
+ comparator_v6_0/CLK io_clamp_low[1] io_clamp_high[1] sky130_fd_sc_hd__buf_16
Xsky130_fd_sc_hd__buf_2_4 io_analog[1] io_clamp_low[1] io_clamp_high[1] sky130_fd_sc_hd__buf_2_4/X
+ io_clamp_low[1] io_clamp_high[1] sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_16_4 sky130_fd_sc_hd__buf_2_4/X io_clamp_low[1] io_clamp_high[1]
+ io_analog[0] io_clamp_low[1] io_clamp_high[1] sky130_fd_sc_hd__buf_16
Xcomparator_v6_0 comparator_v6_0/Outn io_analog[5] io_analog[6] comparator_v6_0/CLK
+ io_clamp_high[1] io_clamp_low[1] comparator_v6_0/Outp comparator_v6_0/CLKBAR comparator_v6
V0 io_clamp_high[1] vccd1 0.0
V1 io_clamp_high[1] io_clamp_high[2] 0.0
V2 io_clamp_low[1] io_clamp_low[2] 0.0
V3 io_clamp_low[1] vssa1 0.0
C0 io_clamp_high[1] sky130_fd_sc_hd__buf_2_1/X 66.21fF
C1 io_clamp_high[1] io_analog[0] 115.74fF
C2 m4_175894_702434# io_analog[6] 48.42fF
C3 m4_180902_677200# io_analog[6] 104.05fF
C4 io_analog[6] m4_165578_698240# 125.98fF
C5 io_clamp_high[1] comparator_v6_0/Outn 9.36fF
C6 sky130_fd_sc_hd__buf_2_3/X m4_204098_586508# 4.77fF
C7 m4_186716_584374# io_analog[6] 185.47fF
C8 io_clamp_high[1] sky130_fd_sc_hd__buf_2_3/X 122.04fF
C9 sky130_fd_sc_hd__buf_2_0/X io_clamp_high[1] 66.26fF
C10 m4_170578_677212# io_analog[6] 53.59fF
C11 io_clamp_high[1] io_analog[3] 34.41fF
C12 io_clamp_high[1] io_analog[6] 111.81fF
C13 m4_204098_586508# io_analog[5] 176.62fF
C14 comparator_v6_0/CLKBAR io_analog[5] 2.23fF
C15 io_clamp_high[1] io_analog[5] 155.94fF
C16 io_clamp_high[1] m4_170578_677212# 30.18fF
C17 sky130_fd_sc_hd__buf_2_3/X m4_186716_584374# 4.20fF
C18 comparator_v6_0/CLK io_analog[6] 2.17fF
C19 sky130_fd_sc_hd__buf_2_3/X io_analog[5] 75.68fF
C20 sky130_fd_sc_hd__buf_2_2/X m4_186716_584374# 4.20fF
C21 io_analog[4] io_clamp_low[1] 25.05fF
C22 vssa1 io_clamp_low[1] 14.37fF
C23 vssd2 io_clamp_low[1] 13.04fF
C24 vssd1 io_clamp_low[1] 13.62fF
C25 vdda2 io_clamp_low[1] 13.04fF
C26 vdda1 io_clamp_low[1] 26.08fF
C27 vssa2 io_clamp_low[1] 13.04fF
C28 vccd2 io_clamp_low[1] 13.04fF
C29 io_analog[10] io_clamp_low[1] 6.83fF
C30 io_clamp_high[0] io_clamp_low[1] 3.58fF
C31 io_clamp_low[0] io_clamp_low[1] 3.58fF
C32 io_analog[9] io_clamp_low[1] 6.83fF
C33 m4_141154_541976# io_clamp_low[1] 136.63fF **FLOATING
C34 m4_204098_586508# io_clamp_low[1] 29.23fF **FLOATING
C35 m4_186716_584374# io_clamp_low[1] 28.89fF **FLOATING
C36 m4_180902_677200# io_clamp_low[1] 18.04fF **FLOATING
C37 m4_170578_677212# io_clamp_low[1] 32.74fF **FLOATING
C38 m4_165578_698240# io_clamp_low[1] 4.28fF **FLOATING
C39 io_analog[3] io_clamp_low[1] 26.43fF
C40 io_clamp_high[1] io_clamp_low[1] 2789.92fF
C41 comparator_v6_0/Outp io_clamp_low[1] 26.62fF
C42 comparator_v6_0/Outn io_clamp_low[1] 19.87fF
C43 comparator_v6_0/CLK io_clamp_low[1] 17.79fF
C44 comparator_v6_0/fp io_clamp_low[1] 2.32fF
C45 comparator_v6_0/fn io_clamp_low[1] 2.31fF
C46 io_analog[5] io_clamp_low[1] 358.90fF
C47 io_analog[6] io_clamp_low[1] 282.38fF
C48 comparator_v6_0/Dp io_clamp_low[1] 3.53fF
C49 comparator_v6_0/Dn io_clamp_low[1] 3.23fF
C50 comparator_v6_0/CLKBAR io_clamp_low[1] 7.21fF
C51 io_analog[0] io_clamp_low[1] 431.97fF
C52 io_analog[1] io_clamp_low[1] 25.06fF
C53 sky130_fd_sc_hd__buf_2_2/X io_clamp_low[1] 354.67fF
C54 io_analog[7] io_clamp_low[1] 64.66fF
C55 sky130_fd_sc_hd__buf_2_3/X io_clamp_low[1] 303.55fF
C56 io_analog[8] io_clamp_low[1] 68.13fF
C57 io_analog[2] io_clamp_low[1] 25.67fF
C58 sky130_fd_sc_hd__buf_2_1/X io_clamp_low[1] 190.70fF
C59 sky130_fd_sc_hd__buf_2_0/X io_clamp_low[1] 195.71fF
.ends

