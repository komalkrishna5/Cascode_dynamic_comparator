magic
tech sky130A
magscale 1 2
timestamp 1651835070
<< nmos >>
rect -63 -450 -33 -350
rect 33 -450 63 -350
<< ndiff >>
rect -121 -361 -63 -350
rect -125 -373 -63 -361
rect -125 -427 -113 -373
rect -79 -427 -63 -373
rect -125 -439 -63 -427
rect -121 -450 -63 -439
rect -33 -373 33 -350
rect -33 -427 -17 -373
rect 17 -427 33 -373
rect -33 -450 33 -427
rect 63 -361 121 -350
rect 63 -373 125 -361
rect 63 -427 79 -373
rect 113 -427 125 -373
rect 63 -439 125 -427
rect 63 -450 121 -439
<< ndiffc >>
rect -113 -427 -79 -373
rect -17 -427 17 -373
rect 79 -427 113 -373
<< poly >>
rect -63 -350 -33 -324
rect 33 -350 63 -324
rect -63 -476 -33 -450
rect 33 -476 63 -450
<< locali >>
rect -113 -373 -79 -357
rect -113 -443 -79 -427
rect -17 -373 17 -357
rect -17 -443 17 -427
rect 79 -373 113 -357
rect 79 -443 113 -427
<< viali >>
rect -113 -427 -79 -373
rect -17 -427 17 -373
rect 79 -427 113 -373
<< metal1 >>
rect -119 -373 -73 -361
rect -119 -427 -113 -373
rect -79 -427 -73 -373
rect -119 -439 -73 -427
rect -23 -373 23 -361
rect -23 -427 -17 -373
rect 17 -427 23 -373
rect -23 -439 23 -427
rect 73 -373 119 -361
rect 73 -427 79 -373
rect 113 -427 119 -373
rect 73 -439 119 -427
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 0.5 l 0.150 m 1 nf 2 diffcov 70 polycov 70 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 70 rlcov 70 topc 1 botc 0 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 0 viasrc 70 viadrn 70 viagate 70 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
