magic
tech sky130A
magscale 1 2
timestamp 1651918812
<< nwell >>
rect -351 74 337 460
rect -161 -356 163 74
<< pmos >>
rect -63 -250 -33 250
rect 33 -250 63 250
<< pdiff >>
rect -125 238 -63 250
rect -125 -238 -113 238
rect -79 -238 -63 238
rect -125 -250 -63 -238
rect -33 238 33 250
rect -33 -238 -17 238
rect 17 -238 33 238
rect -33 -250 33 -238
rect 63 238 125 250
rect 63 -238 79 238
rect 113 -238 125 238
rect 63 -250 125 -238
<< pdiffc >>
rect -113 -238 -79 238
rect -17 -238 17 238
rect 79 -238 113 238
<< poly >>
rect -63 250 -33 276
rect 33 250 63 278
rect -63 -280 -33 -250
rect 33 -276 63 -250
<< locali >>
rect -113 238 -79 254
rect -113 -254 -79 -238
rect -17 238 17 254
rect -17 -254 17 -238
rect 79 238 113 254
rect 79 -254 113 -238
<< viali >>
rect -113 -167 -79 167
rect -17 -167 17 167
rect 79 -167 113 167
<< metal1 >>
rect -119 167 -73 179
rect -119 -167 -113 167
rect -79 -167 -73 167
rect -119 -179 -73 -167
rect -23 167 23 179
rect -23 -167 -17 167
rect 17 -167 23 167
rect -23 -179 23 -167
rect 73 167 119 179
rect 73 -167 79 167
rect 113 -167 119 167
rect 73 -179 119 -167
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 2.5 l 0.15 m 1 nf 2 diffcov 100 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 0 botc 0 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 0 viasrc 70 viadrn 70 viagate 70 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
