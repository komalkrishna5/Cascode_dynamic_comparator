magic
tech sky130A
magscale 1 2
timestamp 1651470485
<< nwell >>
rect -319 -202 169 204
<< pmos >>
rect -63 -100 -33 100
rect 33 -100 63 100
<< pdiff >>
rect -139 62 -63 100
rect -139 -62 -113 62
rect -79 -62 -63 62
rect -139 -100 -63 -62
rect -33 62 33 100
rect -33 -62 -17 62
rect 17 -62 33 62
rect -33 -100 33 -62
rect 63 74 121 100
rect 63 62 125 74
rect 63 -62 79 62
rect 113 -62 125 62
rect 63 -74 125 -62
rect 63 -100 121 -74
<< pdiffc >>
rect -113 -62 -79 62
rect -17 -62 17 62
rect 79 -62 113 62
<< poly >>
rect -63 100 -33 126
rect 33 100 63 126
rect -63 -130 -33 -100
rect 33 -130 63 -100
<< locali >>
rect -139 62 -79 78
rect -139 -62 -113 62
rect -139 -78 -79 -62
rect -17 62 17 78
rect -17 -78 17 -62
rect 79 62 113 78
rect 79 -78 113 -62
<< viali >>
rect -113 -44 -79 44
rect 79 -44 113 44
<< metal1 >>
rect -119 44 -73 56
rect -119 -44 -113 44
rect -79 -44 -73 44
rect -119 -56 -73 -44
rect 73 44 119 56
rect 73 -44 79 44
rect 113 -44 119 44
rect 73 -56 119 -44
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 1 l 0.15 m 1 nf 2 diffcov 70 polycov 70 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 70 rlcov 70 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 0 viasrc 50 viadrn 50 viagate 50 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
