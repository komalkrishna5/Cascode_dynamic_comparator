magic
tech sky130A
magscale 1 2
timestamp 1654411931
use inv_W1#0  inv_W1_0 ~/mycomparator_copy1/layout/myinv_layout2
timestamp 0
transform 1 0 100 0 1 72
box 0 0 1 1
use inv_W2#0  inv_W2_0
timestamp 1647355571
transform 1 0 588 0 1 72
box -120 -72 404 878
<< end >>
