magic
tech sky130A
magscale 1 2
timestamp 1652163895
<< nwell >>
rect -720 994 1018 1328
<< poly >>
rect -462 912 -432 1040
rect -506 870 -432 912
rect 706 910 738 1040
rect 706 862 780 910
rect -168 700 -42 720
rect -168 654 -148 700
rect -72 654 -42 700
rect -168 604 -42 654
rect 316 688 446 714
rect 316 650 338 688
rect 418 650 446 688
rect 316 614 446 650
rect 318 602 348 614
rect 414 588 444 614
rect -168 234 -138 264
rect -72 236 -42 266
rect 318 256 348 264
rect 414 256 444 264
rect -656 -74 -594 -58
rect -656 -116 -640 -74
rect -606 -116 -594 -74
rect -656 -132 -594 -116
rect 864 -72 926 -56
rect 864 -114 880 -72
rect 914 -114 926 -72
rect 864 -130 926 -114
rect -640 -158 -610 -132
rect 882 -166 912 -130
rect -434 -396 -404 -394
rect -338 -396 -308 -394
rect -242 -396 -212 -394
rect -146 -396 -116 -394
rect -434 -568 -116 -396
rect -434 -634 -406 -568
rect -144 -634 -116 -568
rect -434 -660 -116 -634
rect 80 -570 206 -342
rect 80 -638 104 -570
rect 180 -638 206 -570
rect 80 -658 206 -638
rect 388 -402 418 -396
rect 484 -402 514 -396
rect 580 -402 610 -396
rect 676 -402 706 -396
rect 388 -564 706 -402
rect 388 -634 414 -564
rect 680 -634 706 -564
rect 388 -660 706 -634
<< polycont >>
rect -148 654 -72 700
rect 338 650 418 688
rect -640 -116 -606 -74
rect 880 -114 914 -72
rect -406 -634 -144 -568
rect 104 -638 180 -570
rect 414 -634 680 -564
<< locali >>
rect -720 1336 1020 1386
rect -508 1208 -474 1336
rect 748 1210 782 1336
rect 314 820 442 832
rect 314 782 330 820
rect 426 782 442 820
rect -164 708 -56 716
rect -164 644 -158 708
rect -60 644 -56 708
rect -164 638 -56 644
rect 314 714 442 782
rect 314 688 446 714
rect 314 650 338 688
rect 418 650 446 688
rect 314 636 446 650
rect 316 634 446 636
rect -218 234 -184 548
rect -26 234 8 546
rect 92 234 182 242
rect 268 234 302 280
rect 460 234 494 296
rect -218 230 494 234
rect -218 192 104 230
rect 92 190 104 192
rect 172 192 494 230
rect 172 190 182 192
rect 92 180 182 190
rect -656 -74 -594 -58
rect -656 -116 -642 -74
rect -606 -116 -594 -74
rect -656 -132 -594 -116
rect 864 -72 926 -56
rect 864 -114 878 -72
rect 914 -114 926 -72
rect -484 -162 -66 -128
rect -718 -356 -652 -200
rect -484 -212 -450 -162
rect -292 -206 -258 -162
rect -100 -210 -66 -162
rect 338 -162 756 -128
rect 864 -130 926 -114
rect 338 -208 372 -162
rect 530 -206 564 -162
rect 722 -208 756 -162
rect -598 -422 -564 -348
rect 30 -352 66 -312
rect 122 -313 166 -252
rect 222 -352 256 -314
rect 30 -422 256 -352
rect 836 -422 870 -346
rect 954 -358 1020 -202
rect -720 -474 1020 -422
rect -422 -566 -128 -550
rect -422 -634 -406 -566
rect -144 -634 -128 -566
rect -422 -652 -128 -634
rect 78 -570 206 -552
rect 78 -638 104 -570
rect 180 -638 206 -570
rect 78 -660 206 -638
rect 398 -564 696 -548
rect 398 -634 414 -564
rect 680 -634 696 -564
rect 398 -650 696 -634
<< viali >>
rect 330 782 426 820
rect -158 700 -60 708
rect -158 654 -148 700
rect -148 654 -72 700
rect -72 654 -60 700
rect -158 644 -60 654
rect 104 190 172 230
rect -642 -116 -640 -74
rect -640 -116 -606 -74
rect 878 -114 880 -72
rect 880 -114 914 -72
rect -406 -568 -144 -566
rect -406 -634 -144 -568
rect 106 -638 180 -570
rect 414 -634 680 -564
<< metal1 >>
rect -428 830 -380 1104
rect 314 830 442 832
rect -428 820 442 830
rect -428 810 330 820
rect -430 782 330 810
rect 426 782 442 820
rect -656 -74 -594 -58
rect -430 -70 -380 782
rect 314 770 442 782
rect -168 708 -46 722
rect -168 644 -158 708
rect -60 698 -46 708
rect 654 698 702 1132
rect -60 650 702 698
rect -60 644 -46 650
rect -168 630 -46 644
rect -430 -74 -160 -70
rect -718 -116 -642 -74
rect -606 -116 -160 -74
rect -656 -132 -594 -116
rect -692 -210 -648 -188
rect -390 -246 -352 -116
rect -198 -250 -160 -116
rect -122 -128 -88 468
rect 88 230 194 250
rect 88 190 104 230
rect 172 190 194 230
rect 88 172 194 190
rect -128 -164 -66 -128
rect -104 -262 -66 -164
rect 120 -284 166 172
rect 364 -128 398 350
rect 654 -74 702 650
rect 864 -72 926 -56
rect 864 -74 878 -72
rect 434 -114 878 -74
rect 914 -74 926 -72
rect 914 -114 1020 -74
rect 434 -116 1020 -114
rect 338 -162 406 -128
rect 338 -220 374 -162
rect 434 -212 470 -116
rect 624 -208 660 -116
rect 864 -130 926 -116
rect -422 -566 -128 -550
rect -422 -634 -406 -566
rect -144 -634 -128 -566
rect -422 -654 -128 -634
rect 78 -570 206 -552
rect 78 -638 106 -570
rect 180 -638 206 -570
rect 78 -658 206 -638
rect 398 -564 696 -548
rect 398 -634 414 -564
rect 680 -634 696 -564
rect 398 -650 696 -634
use sky130_fd_pr__nfet_01v8_8FHE5N  sky130_fd_pr__nfet_01v8_8FHE5N_0
timestamp 1651835070
transform 1 0 143 0 1 126
box -125 -476 125 -324
use sky130_fd_pr__nfet_01v8_F5U58G#1  sky130_fd_pr__nfet_01v8_F5U58G_0
timestamp 1651835070
transform 1 0 -625 0 1 116
box -73 -526 73 -274
use sky130_fd_pr__nfet_01v8_F5U58G#1  sky130_fd_pr__nfet_01v8_F5U58G_1
timestamp 1651835070
transform 1 0 897 0 1 120
box -73 -526 73 -274
use sky130_fd_pr__nfet_01v8_G6PLX8  sky130_fd_pr__nfet_01v8_G6PLX8_0
timestamp 1651835070
transform 1 0 -275 0 1 122
box -221 -526 221 -250
use sky130_fd_pr__nfet_01v8_G6PLX8  sky130_fd_pr__nfet_01v8_G6PLX8_1
timestamp 1651835070
transform 1 0 547 0 1 122
box -221 -526 221 -250
use sky130_fd_pr__nfet_01v8_RURP52  sky130_fd_pr__nfet_01v8_RURP52_0
timestamp 1651837652
transform 1 0 -105 0 1 630
box -125 -374 125 -22
use sky130_fd_pr__nfet_01v8_RURP52  sky130_fd_pr__nfet_01v8_RURP52_1
timestamp 1651837652
transform 1 0 381 0 1 630
box -125 -374 125 -22
use sky130_fd_pr__pfet_01v8_RFM3CD#0  sky130_fd_pr__pfet_01v8_RFM3CD_0
timestamp 1646431323
transform 1 0 -447 0 1 1160
box -109 -162 109 162
use sky130_fd_pr__pfet_01v8_RFM3CD#0  sky130_fd_pr__pfet_01v8_RFM3CD_1
timestamp 1646431323
transform 1 0 721 0 1 1160
box -109 -162 109 162
<< end >>
