magic
tech sky130A
magscale 1 2
timestamp 1653304099
<< error_p >>
rect 48 48 78 54
use sky130_fd_pr__nfet_01v8_7RYEVP  sky130_fd_pr__nfet_01v8_7RYEVP_0 ~/my_sky130_project/mag/myinv_layout2
timestamp 1651470485
transform 1 0 63 0 1 143
box -73 -95 73 157
<< end >>
