magic
tech sky130A
magscale 1 2
timestamp 1652082874
<< error_p >>
rect -247 136 -137 162
rect -247 130 297 136
rect 305 130 465 162
rect -269 94 269 100
rect -439 -128 -305 40
rect -271 -198 299 56
rect 305 -198 467 40
<< nwell >>
rect -305 130 -247 162
rect 297 130 305 162
rect -305 -128 305 130
rect -305 -198 -271 -128
rect 299 -198 305 -128
rect -305 -200 305 -198
<< pmos >>
rect -207 -100 -177 100
rect -111 -100 -81 100
rect -15 -100 15 100
rect 81 -100 111 100
rect 177 -100 207 100
<< pdiff >>
rect -269 88 -207 100
rect -269 -88 -257 88
rect -223 -88 -207 88
rect -269 -100 -207 -88
rect -177 88 -111 100
rect -177 -88 -161 88
rect -127 -88 -111 88
rect -177 -100 -111 -88
rect -81 88 -15 100
rect -81 -88 -65 88
rect -31 -88 -15 88
rect -81 -100 -15 -88
rect 15 88 81 100
rect 15 -88 31 88
rect 65 -88 81 88
rect 15 -100 81 -88
rect 111 88 177 100
rect 111 -88 127 88
rect 161 -88 177 88
rect 111 -100 177 -88
rect 207 88 269 100
rect 207 -88 223 88
rect 257 -88 269 88
rect 207 -100 269 -88
<< pdiffc >>
rect -257 -88 -223 88
rect -161 -88 -127 88
rect -65 -88 -31 88
rect 31 -88 65 88
rect 127 -88 161 88
rect 223 -88 257 88
<< poly >>
rect -207 100 -177 126
rect -111 100 -81 130
rect -15 100 15 126
rect 81 100 111 130
rect 177 100 207 126
rect -207 -128 -177 -100
rect -111 -126 -81 -100
rect -15 -128 15 -100
rect 81 -126 111 -100
rect 177 -128 207 -100
<< locali >>
rect -257 88 -223 104
rect -257 -104 -223 -88
rect -161 88 -127 104
rect -161 -104 -127 -88
rect -65 88 -31 104
rect -65 -104 -31 -88
rect 31 88 65 104
rect 31 -104 65 -88
rect 127 88 161 104
rect 127 -104 161 -88
rect 223 88 257 104
rect 223 -104 257 -88
<< viali >>
rect -257 -62 -223 62
rect -161 -62 -127 62
rect -65 -62 -31 62
rect 31 -62 65 62
rect 127 -62 161 62
rect 223 -62 257 62
<< metal1 >>
rect -263 62 -217 74
rect -263 -62 -257 62
rect -223 -62 -217 62
rect -263 -74 -217 -62
rect -167 62 -121 74
rect -167 -62 -161 62
rect -127 -62 -121 62
rect -167 -74 -121 -62
rect -71 62 -25 74
rect -71 -62 -65 62
rect -31 -62 -25 62
rect -71 -74 -25 -62
rect 25 62 71 74
rect 25 -62 31 62
rect 65 -62 71 62
rect 25 -74 71 -62
rect 121 62 167 74
rect 121 -62 127 62
rect 161 -62 167 62
rect 121 -74 167 -62
rect 217 62 263 74
rect 217 -62 223 62
rect 257 -62 263 62
rect 217 -74 263 -62
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 1 l 0.15 m 1 nf 5 diffcov 100 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 0 botc 0 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 0 viasrc 70 viadrn 70 viagate 70 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
