magic
tech sky130A
magscale 1 2
timestamp 1651835070
<< error_p >>
rect -159 -526 -129 -522
rect -63 -526 -33 -522
rect 33 -526 63 -522
rect 129 -526 159 -522
<< nmos >>
rect -159 -500 -129 -300
rect -63 -500 -33 -300
rect 33 -500 63 -300
rect 129 -500 159 -300
<< ndiff >>
rect -217 -326 -159 -300
rect -221 -338 -159 -326
rect -221 -462 -209 -338
rect -175 -462 -159 -338
rect -221 -474 -159 -462
rect -217 -500 -159 -474
rect -129 -338 -63 -300
rect -129 -462 -113 -338
rect -79 -462 -63 -338
rect -129 -500 -63 -462
rect -33 -338 33 -300
rect -33 -462 -17 -338
rect 17 -462 33 -338
rect -33 -500 33 -462
rect 63 -338 129 -300
rect 63 -462 79 -338
rect 113 -462 129 -338
rect 63 -500 129 -462
rect 159 -326 217 -300
rect 159 -338 221 -326
rect 159 -462 175 -338
rect 209 -462 221 -338
rect 159 -474 221 -462
rect 159 -500 217 -474
<< ndiffc >>
rect -209 -462 -175 -338
rect -113 -462 -79 -338
rect -17 -462 17 -338
rect 79 -462 113 -338
rect 175 -462 209 -338
<< poly >>
rect -159 -280 159 -250
rect -159 -300 -129 -280
rect -63 -300 -33 -280
rect 33 -300 63 -280
rect 129 -300 159 -280
rect -159 -522 -129 -500
rect -63 -522 -33 -500
rect 33 -522 63 -500
rect 129 -522 159 -500
<< locali >>
rect -209 -338 -175 -322
rect -209 -478 -175 -462
rect -113 -338 -79 -322
rect -113 -478 -79 -462
rect -17 -338 17 -322
rect -17 -478 17 -462
rect 79 -338 113 -322
rect 79 -478 113 -462
rect 175 -338 209 -322
rect 175 -478 209 -462
<< viali >>
rect -209 -462 -175 -338
rect -113 -462 -79 -338
rect -17 -462 17 -338
rect 79 -462 113 -338
rect 175 -462 209 -338
<< metal1 >>
rect -215 -338 -169 -326
rect -215 -462 -209 -338
rect -175 -462 -169 -338
rect -215 -474 -169 -462
rect -119 -338 -73 -326
rect -119 -462 -113 -338
rect -79 -462 -73 -338
rect -119 -474 -73 -462
rect -23 -338 23 -326
rect -23 -462 -17 -338
rect 17 -462 23 -338
rect -23 -474 23 -462
rect 73 -338 119 -326
rect 73 -462 79 -338
rect 113 -462 119 -338
rect 73 -474 119 -462
rect 169 -338 215 -326
rect 169 -462 175 -338
rect 209 -462 215 -338
rect 169 -474 215 -462
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 1 l 0.150 m 1 nf 4 diffcov 70 polycov 70 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 70 rlcov 70 topc 0 botc 0 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 0 viasrc 70 viadrn 70 viagate 70 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
