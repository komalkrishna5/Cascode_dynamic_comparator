magic
tech sky130A
magscale 1 2
timestamp 1654429859
<< nwell >>
rect 415156 686850 415500 686862
rect 415156 686674 415504 686850
rect 467114 686536 467436 686824
rect 440076 655268 440396 655476
rect 448734 655462 448948 655486
rect 448660 655336 448980 655462
rect 135002 599506 136140 599832
rect 86264 585822 87030 585824
rect 86014 585502 87030 585822
rect 86014 585500 86274 585502
rect 103604 567702 103892 568026
rect 110034 567782 110676 568118
<< nsubdiff >>
rect 415238 686750 415262 686804
rect 415362 686750 415386 686804
rect 467192 686674 467216 686726
rect 467330 686674 467354 686726
rect 440186 655360 440210 655420
rect 440320 655360 440344 655420
rect 448760 655394 448784 655432
rect 448874 655394 448898 655432
rect 135308 599714 135352 599738
rect 135308 599572 135352 599596
rect 86102 585728 86156 585752
rect 86102 585592 86156 585616
rect 110358 568032 110426 568056
rect 103728 567908 103784 567932
rect 110358 567876 110426 567900
rect 103728 567782 103784 567806
<< nsubdiffcont >>
rect 415262 686750 415362 686804
rect 467216 686674 467330 686726
rect 440210 655360 440320 655420
rect 448784 655394 448874 655432
rect 135308 599596 135352 599714
rect 86102 585616 86156 585728
rect 103728 567806 103784 567908
rect 110358 567900 110426 568032
<< locali >>
rect 467316 691416 467882 691454
rect 415478 691358 415536 691360
rect 415416 691316 415982 691358
rect 415416 691208 415460 691316
rect 415562 691208 415820 691316
rect 415922 691208 415982 691316
rect 415416 691076 415982 691208
rect 415416 690968 415460 691076
rect 415562 690968 415820 691076
rect 415922 690968 415982 691076
rect 467316 691308 467360 691416
rect 467462 691308 467720 691416
rect 467822 691308 467882 691416
rect 467316 691176 467882 691308
rect 467316 691068 467360 691176
rect 467462 691068 467720 691176
rect 467822 691068 467882 691176
rect 467316 691026 467882 691068
rect 415416 690926 415982 690968
rect 415476 690760 415534 690926
rect 415434 688844 415560 690760
rect 467430 690536 467494 691026
rect 467420 690510 467494 690536
rect 467420 688806 467492 690510
rect 412670 688608 414760 688612
rect 412670 688376 415206 688608
rect 465730 688604 466792 688608
rect 412670 688212 413812 688376
rect 413996 688212 414212 688376
rect 414394 688212 415206 688376
rect 412670 687976 415206 688212
rect 412670 687812 413812 687976
rect 413996 687812 414212 687976
rect 414394 687812 415206 687976
rect 412670 687576 415206 687812
rect 412670 687412 413812 687576
rect 413996 687412 414212 687576
rect 414394 687412 415206 687576
rect 412670 687176 415206 687412
rect 412670 687012 413812 687176
rect 413996 687012 414212 687176
rect 414394 687012 415206 687176
rect 412670 686948 415206 687012
rect 412670 686942 414760 686948
rect 414930 686946 415206 686948
rect 415774 688586 416000 688592
rect 416130 688586 416872 688598
rect 415774 688376 416872 688586
rect 415774 688212 416212 688376
rect 416396 688212 416612 688376
rect 416796 688212 416872 688376
rect 415774 687976 416872 688212
rect 415774 687812 416212 687976
rect 416396 687812 416612 687976
rect 416796 687812 416872 687976
rect 415774 687576 416872 687812
rect 415774 687412 416212 687576
rect 416396 687412 416612 687576
rect 416796 687412 416872 687576
rect 415774 687176 416872 687412
rect 415774 687012 416212 687176
rect 416396 687012 416622 687176
rect 416806 687012 416872 687176
rect 415330 686868 415404 686946
rect 415774 686944 416872 687012
rect 465730 688376 467146 688604
rect 465730 688212 465812 688376
rect 465996 688212 466212 688376
rect 466370 688212 467146 688376
rect 465730 687976 467146 688212
rect 465730 687812 465812 687976
rect 465996 687812 466212 687976
rect 466370 687812 467146 687976
rect 465730 687576 467146 687812
rect 465730 687412 465812 687576
rect 465996 687412 466212 687576
rect 466370 687412 467146 687576
rect 465730 687176 467146 687412
rect 465730 687012 465812 687176
rect 465996 687012 466212 687176
rect 466370 687012 467146 687176
rect 465730 686948 467146 687012
rect 467712 688586 468086 688592
rect 468130 688586 468872 688598
rect 467712 688376 468872 688586
rect 467712 688212 468212 688376
rect 468396 688212 468612 688376
rect 468796 688212 468872 688376
rect 467712 687976 468872 688212
rect 467712 687812 468212 687976
rect 468396 687812 468612 687976
rect 468796 687812 468872 687976
rect 467712 687576 468872 687812
rect 467712 687412 468212 687576
rect 468396 687412 468612 687576
rect 468796 687412 468872 687576
rect 467712 687176 468872 687412
rect 467712 687012 468212 687176
rect 468396 687012 468622 687176
rect 468806 687012 468872 687176
rect 465730 686944 466598 686948
rect 467712 686944 468872 687012
rect 415774 686936 416238 686944
rect 467712 686936 468238 686944
rect 415300 686804 415406 686868
rect 415246 686750 415262 686804
rect 415362 686750 415406 686804
rect 415300 686748 415406 686750
rect 415508 686508 415546 686926
rect 415774 686924 416000 686936
rect 467712 686928 468086 686936
rect 467268 686726 467332 686888
rect 467200 686674 467216 686726
rect 467330 686674 467346 686726
rect 467268 686672 467332 686674
rect 415502 686258 415546 686508
rect 415502 685916 415540 686258
rect 467442 686018 467478 686872
rect 467440 685926 467478 686018
rect 415494 685558 415552 685916
rect 467440 685732 467476 685926
rect 467364 685590 467548 685732
rect 415416 685516 415982 685558
rect 467364 685554 467550 685590
rect 415416 685408 415460 685516
rect 415562 685408 415820 685516
rect 415922 685408 415982 685516
rect 415416 685276 415982 685408
rect 415416 685168 415460 685276
rect 415562 685168 415820 685276
rect 415922 685168 415982 685276
rect 415416 685126 415982 685168
rect 467316 685512 467882 685554
rect 467316 685404 467360 685512
rect 467462 685404 467720 685512
rect 467822 685404 467882 685512
rect 467316 685272 467882 685404
rect 467316 685164 467360 685272
rect 467462 685164 467720 685272
rect 467822 685164 467882 685272
rect 467316 685122 467882 685164
rect 440216 657716 440782 657758
rect 440216 657608 440260 657716
rect 440362 657608 440620 657716
rect 440722 657608 440782 657716
rect 440216 657476 440782 657608
rect 440216 657368 440260 657476
rect 440362 657368 440620 657476
rect 440722 657368 440782 657476
rect 440216 657328 440782 657368
rect 448816 657716 449382 657758
rect 448816 657608 448860 657716
rect 448962 657608 449220 657716
rect 449322 657608 449382 657716
rect 448816 657476 449382 657608
rect 448816 657368 448860 657476
rect 448962 657368 449220 657476
rect 449322 657368 449382 657476
rect 448816 657328 449382 657368
rect 437730 656602 438598 656608
rect 437730 656600 439968 656602
rect 437730 656376 440108 656600
rect 437730 656212 437812 656376
rect 437996 656212 438212 656376
rect 438396 656212 440108 656376
rect 437730 655976 440108 656212
rect 440372 656150 440470 657328
rect 448972 657212 449070 657328
rect 442330 656700 443072 656712
rect 442232 656490 443072 656700
rect 442232 656326 442412 656490
rect 442596 656326 442812 656490
rect 442996 656326 443072 656490
rect 440640 656184 441194 656190
rect 442232 656184 443072 656326
rect 437730 655812 437812 655976
rect 437996 655812 438212 655976
rect 438396 655812 440108 655976
rect 437730 655576 440108 655812
rect 440398 655746 440434 656150
rect 440640 656090 443072 656184
rect 440640 655926 442412 656090
rect 442596 655926 442812 656090
rect 442996 655926 443072 656090
rect 437730 655412 437812 655576
rect 437996 655412 438212 655576
rect 438396 655420 440108 655576
rect 440640 655690 443072 655926
rect 438396 655412 440210 655420
rect 437730 655362 440210 655412
rect 437730 655176 440108 655362
rect 440194 655360 440210 655362
rect 440320 655360 440336 655420
rect 440396 655236 440446 655544
rect 440640 655526 442412 655690
rect 442596 655526 442812 655690
rect 442996 655526 443072 655690
rect 440640 655290 443072 655526
rect 437730 655012 437812 655176
rect 437996 655012 438212 655176
rect 438396 655012 440108 655176
rect 440394 655080 440450 655236
rect 440640 655196 442412 655290
rect 440640 655192 441194 655196
rect 442232 655126 442412 655196
rect 442596 655126 442822 655290
rect 443006 655126 443072 655290
rect 437730 654944 440108 655012
rect 438466 654934 440108 654944
rect 439784 654930 440108 654934
rect 440368 654758 440486 655080
rect 442232 655058 443072 655126
rect 446130 656602 446998 656608
rect 446130 656376 448714 656602
rect 446130 656212 446212 656376
rect 446396 656212 446612 656376
rect 446796 656212 448714 656376
rect 446130 655976 448714 656212
rect 448972 656176 449072 657212
rect 450730 656700 451472 656712
rect 450632 656490 451472 656700
rect 450632 656326 450812 656490
rect 450996 656326 451212 656490
rect 451396 656326 451472 656490
rect 450632 656184 451472 656326
rect 450628 656180 451472 656184
rect 446130 655812 446212 655976
rect 446396 655812 446612 655976
rect 446796 655812 448714 655976
rect 446130 655576 448714 655812
rect 448986 655746 449022 656176
rect 449226 656090 451472 656180
rect 449226 655926 450814 656090
rect 450996 655926 451212 656090
rect 451396 655926 451472 656090
rect 446130 655412 446212 655576
rect 446396 655412 446612 655576
rect 446796 655440 448714 655576
rect 449226 655690 451472 655926
rect 449226 655526 450814 655690
rect 450996 655526 451212 655690
rect 451396 655526 451472 655690
rect 446796 655432 448818 655440
rect 446796 655412 448784 655432
rect 446130 655394 448784 655412
rect 448874 655394 448890 655432
rect 446130 655382 448818 655394
rect 446130 655176 448714 655382
rect 448972 655210 449046 655514
rect 449226 655290 451472 655526
rect 442232 655050 442438 655058
rect 446130 655012 446212 655176
rect 446396 655012 446612 655176
rect 446796 655012 448714 655176
rect 446130 654944 448714 655012
rect 446866 654934 448714 654944
rect 447078 654924 448714 654934
rect 448966 654876 449086 655210
rect 449226 655190 450814 655290
rect 449226 655184 449590 655190
rect 450632 655126 450812 655190
rect 450996 655126 451222 655290
rect 451406 655126 451472 655290
rect 450632 655058 451472 655126
rect 450632 655050 450838 655058
rect 448968 654758 449086 654876
rect 440216 654716 440782 654758
rect 440216 654608 440260 654716
rect 440362 654608 440620 654716
rect 440722 654608 440782 654716
rect 440216 654476 440782 654608
rect 440216 654368 440260 654476
rect 440362 654368 440620 654476
rect 440722 654368 440782 654476
rect 440216 654328 440782 654368
rect 448816 654716 449382 654758
rect 448816 654608 448860 654716
rect 448962 654608 449220 654716
rect 449322 654608 449382 654716
rect 448816 654476 449382 654608
rect 448816 654368 448860 654476
rect 448962 654368 449220 654476
rect 449322 654368 449382 654476
rect 448816 654328 449382 654368
rect 134396 600374 139074 600454
rect 134212 600344 139074 600374
rect 134212 600104 134560 600344
rect 134868 600104 135160 600344
rect 135468 600104 135760 600344
rect 136068 600104 136360 600344
rect 136668 600104 136960 600344
rect 137268 600104 137560 600344
rect 137868 600104 138160 600344
rect 138468 600104 139074 600344
rect 134212 599978 139074 600104
rect 134212 599972 139038 599978
rect 135308 599730 135350 599972
rect 135308 599714 135352 599730
rect 133984 599596 134258 599606
rect 133984 599540 134006 599596
rect 134086 599540 134126 599596
rect 134206 599540 134258 599596
rect 135308 599580 135352 599596
rect 140384 599596 140628 599606
rect 133984 599510 134258 599540
rect 138120 599550 139236 599556
rect 138120 599544 140298 599550
rect 140384 599546 140406 599596
rect 140370 599544 140406 599546
rect 138120 599540 140406 599544
rect 140486 599540 140526 599596
rect 140606 599540 140628 599596
rect 133984 599496 134664 599510
rect 133984 599440 134006 599496
rect 134086 599440 134126 599496
rect 134206 599442 134664 599496
rect 134864 599468 136198 599502
rect 138120 599496 140628 599540
rect 138120 599488 140406 599496
rect 138120 599478 140298 599488
rect 138120 599476 139236 599478
rect 134206 599440 134258 599442
rect 133984 599410 134258 599440
rect 140384 599440 140406 599488
rect 140486 599440 140526 599496
rect 140606 599440 140628 599496
rect 140384 599410 140628 599440
rect 134242 599060 134360 599078
rect 134242 599030 139086 599060
rect 134242 598866 134398 599030
rect 134592 598866 134798 599030
rect 134992 598866 135198 599030
rect 135392 598866 135598 599030
rect 135792 598866 135998 599030
rect 136192 598866 136398 599030
rect 136592 598866 136798 599030
rect 136992 598866 137198 599030
rect 137392 598866 137598 599030
rect 137792 598866 137998 599030
rect 138192 598866 138398 599030
rect 138592 598866 138798 599030
rect 138992 598866 139086 599030
rect 134242 598790 139086 598866
rect 134242 598626 134398 598790
rect 134592 598626 134798 598790
rect 134992 598626 135198 598790
rect 135392 598626 135598 598790
rect 135792 598626 135998 598790
rect 136192 598626 136398 598790
rect 136592 598626 136798 598790
rect 136992 598626 137198 598790
rect 137392 598626 137598 598790
rect 137792 598626 137998 598790
rect 138192 598626 138398 598790
rect 138592 598626 138798 598790
rect 138992 598626 139086 598790
rect 134242 598562 139086 598626
rect 85396 586374 90074 586454
rect 85212 586344 90074 586374
rect 85212 586104 85560 586344
rect 85868 586104 86160 586344
rect 86468 586104 86760 586344
rect 87068 586104 87360 586344
rect 87668 586104 87960 586344
rect 88268 586104 88560 586344
rect 88868 586104 89160 586344
rect 89468 586104 90074 586344
rect 85212 585978 90074 586104
rect 424124 586416 424202 586450
rect 424124 586174 424142 586416
rect 424184 586174 424202 586416
rect 85212 585972 90038 585978
rect 424124 585892 424202 586174
rect 85982 585766 86156 585802
rect 86102 585728 86156 585766
rect 84984 585596 85258 585606
rect 86102 585600 86156 585616
rect 84984 585540 85006 585596
rect 85086 585540 85126 585596
rect 85206 585540 85258 585596
rect 91384 585596 91628 585606
rect 84984 585510 85258 585540
rect 89012 585544 91298 585550
rect 91384 585546 91406 585596
rect 91370 585544 91406 585546
rect 89012 585540 91406 585544
rect 91486 585540 91526 585596
rect 91606 585540 91628 585596
rect 84984 585496 85718 585510
rect 84984 585440 85006 585496
rect 85086 585440 85126 585496
rect 85206 585442 85718 585496
rect 85872 585498 86980 585500
rect 85872 585464 87088 585498
rect 89012 585496 91628 585540
rect 89012 585488 91406 585496
rect 89012 585478 91298 585488
rect 89012 585476 90236 585478
rect 85872 585458 85894 585464
rect 86026 585460 87088 585464
rect 86026 585458 86980 585460
rect 85206 585440 85258 585442
rect 84984 585410 85258 585440
rect 91384 585440 91406 585488
rect 91486 585440 91526 585496
rect 91606 585440 91628 585496
rect 91384 585410 91628 585440
rect 85242 585030 90086 585078
rect 85242 584866 85398 585030
rect 85592 584866 85798 585030
rect 85992 584866 86198 585030
rect 86392 584866 86598 585030
rect 86792 584866 86998 585030
rect 87192 584866 87398 585030
rect 87592 584866 87798 585030
rect 87992 584866 88198 585030
rect 88392 584866 88598 585030
rect 88792 584866 88998 585030
rect 89192 584866 89398 585030
rect 89592 584866 89798 585030
rect 89992 584866 90086 585030
rect 85242 584790 90086 584866
rect 424114 585046 424188 585350
rect 424114 584824 424132 585046
rect 424174 584824 424188 585046
rect 424114 584792 424188 584824
rect 85242 584626 85398 584790
rect 85592 584626 85798 584790
rect 85992 584626 86198 584790
rect 86392 584626 86598 584790
rect 86792 584626 86998 584790
rect 87192 584626 87398 584790
rect 87592 584626 87798 584790
rect 87992 584626 88198 584790
rect 88392 584626 88598 584790
rect 88792 584626 88998 584790
rect 89192 584626 89398 584790
rect 89592 584626 89798 584790
rect 89992 584626 90086 584790
rect 85242 584562 90086 584626
rect 101690 568824 106034 568854
rect 107396 568824 111740 568854
rect 101608 568744 106034 568824
rect 101608 568504 101854 568744
rect 102162 568504 102454 568744
rect 102762 568504 103054 568744
rect 103362 568504 103654 568744
rect 103962 568504 104254 568744
rect 104562 568504 104854 568744
rect 105162 568504 105454 568744
rect 105762 568504 106034 568744
rect 101608 568356 106034 568504
rect 101606 568328 106034 568356
rect 107314 568744 111740 568824
rect 107314 568504 107560 568744
rect 107868 568504 108160 568744
rect 108468 568504 108760 568744
rect 109068 568504 109360 568744
rect 109668 568504 109960 568744
rect 110268 568504 110560 568744
rect 110868 568504 111160 568744
rect 111468 568504 111740 568744
rect 101606 568136 106030 568328
rect 107314 568264 111740 568504
rect 107314 568226 111976 568264
rect 103014 567988 104254 568136
rect 108020 568064 110046 568226
rect 110358 568032 110428 568226
rect 103580 567974 103782 567988
rect 103610 567972 103782 567974
rect 103728 567924 103782 567972
rect 103728 567908 103784 567924
rect 110426 567900 110428 568032
rect 110358 567884 110426 567900
rect 113384 567844 113620 567854
rect 102842 567796 103076 567806
rect 102842 567740 102864 567796
rect 102944 567740 102984 567796
rect 103064 567740 103076 567796
rect 103728 567790 103784 567806
rect 103986 567796 104220 567806
rect 102842 567712 103076 567740
rect 103986 567740 104006 567796
rect 104086 567740 104126 567796
rect 104206 567740 104220 567796
rect 103214 567712 103288 567714
rect 102842 567696 103288 567712
rect 103986 567708 104220 567740
rect 103648 567698 104220 567708
rect 102842 567640 102864 567696
rect 102944 567640 102984 567696
rect 103064 567644 103288 567696
rect 103479 567696 104220 567698
rect 103479 567664 104006 567696
rect 103648 567652 104006 567664
rect 103064 567640 103076 567644
rect 102842 567610 103076 567640
rect 103986 567640 104006 567652
rect 104086 567640 104126 567696
rect 104206 567640 104220 567696
rect 103986 567610 104220 567640
rect 106984 567796 107220 567806
rect 106984 567740 107006 567796
rect 107086 567740 107126 567796
rect 107206 567794 107220 567796
rect 109970 567794 113340 567798
rect 113384 567794 113406 567844
rect 107206 567782 107290 567794
rect 109970 567788 113406 567794
rect 113486 567788 113526 567844
rect 113606 567842 113620 567844
rect 113606 567788 113622 567842
rect 109970 567786 113622 567788
rect 107206 567780 107948 567782
rect 107206 567742 108046 567780
rect 109970 567750 113620 567786
rect 113090 567744 113620 567750
rect 107206 567740 107976 567742
rect 106984 567738 107290 567740
rect 113090 567738 113406 567744
rect 106984 567696 107220 567738
rect 106984 567640 107006 567696
rect 107086 567640 107126 567696
rect 107206 567640 107220 567696
rect 113384 567688 113406 567738
rect 113486 567688 113526 567744
rect 113606 567688 113620 567744
rect 113384 567658 113620 567688
rect 106984 567610 107220 567640
rect 107908 567334 110066 567538
rect 101238 567068 106104 567240
rect 101238 566904 101408 567068
rect 101602 566904 101808 567068
rect 102002 566904 102208 567068
rect 102402 566904 102608 567068
rect 102802 566904 103008 567068
rect 103202 566904 103408 567068
rect 103602 566904 103808 567068
rect 104002 566904 104208 567068
rect 104402 566904 104608 567068
rect 104802 566904 105008 567068
rect 105202 566904 105408 567068
rect 105602 566904 105808 567068
rect 106002 566904 106104 567068
rect 101238 566828 106104 566904
rect 101238 566664 101408 566828
rect 101602 566664 101808 566828
rect 102002 566664 102208 566828
rect 102402 566664 102608 566828
rect 102802 566664 103008 566828
rect 103202 566664 103408 566828
rect 103602 566664 103808 566828
rect 104002 566664 104208 566828
rect 104402 566664 104608 566828
rect 104802 566664 105008 566828
rect 105202 566664 105408 566828
rect 105602 566664 105808 566828
rect 106002 566664 106104 566828
rect 101238 566568 106104 566664
rect 107228 567030 112094 567334
rect 107228 566866 107398 567030
rect 107592 566866 107798 567030
rect 107908 567024 110198 567030
rect 107992 566866 108198 567024
rect 108392 566866 108598 567024
rect 108792 566866 108998 567024
rect 109192 566866 109398 567024
rect 109592 566866 109798 567024
rect 109992 566866 110198 567024
rect 110392 566866 110598 567030
rect 110792 566866 110998 567030
rect 111192 566866 111398 567030
rect 111592 566866 111798 567030
rect 111992 566866 112094 567030
rect 107228 566790 112094 566866
rect 107228 566626 107398 566790
rect 107592 566626 107798 566790
rect 107992 566626 108198 566790
rect 108392 566626 108598 566790
rect 108792 566626 108998 566790
rect 109192 566626 109398 566790
rect 109592 566626 109798 566790
rect 109992 566626 110198 566790
rect 110392 566626 110598 566790
rect 110792 566626 110998 566790
rect 111192 566626 111398 566790
rect 111592 566626 111798 566790
rect 111992 566626 112094 566790
rect 107228 566530 112094 566626
<< viali >>
rect 118843 695007 118877 695109
rect 126213 694803 126247 694905
rect 415460 691208 415562 691316
rect 415820 691208 415922 691316
rect 415460 690968 415562 691076
rect 415820 690968 415922 691076
rect 467360 691308 467462 691416
rect 467720 691308 467822 691416
rect 467360 691068 467462 691176
rect 467720 691068 467822 691176
rect 413812 688212 413996 688376
rect 414212 688212 414394 688376
rect 413812 687812 413996 687976
rect 414212 687812 414394 687976
rect 413812 687412 413996 687576
rect 414212 687412 414394 687576
rect 413812 687012 413996 687176
rect 414212 687012 414394 687176
rect 416212 688212 416396 688376
rect 416612 688212 416796 688376
rect 416212 687812 416396 687976
rect 416612 687812 416796 687976
rect 416212 687412 416396 687576
rect 416612 687412 416796 687576
rect 416212 687012 416396 687176
rect 416622 687012 416806 687176
rect 465812 688212 465996 688376
rect 466212 688212 466370 688376
rect 465812 687812 465996 687976
rect 466212 687812 466370 687976
rect 465812 687412 465996 687576
rect 466212 687412 466370 687576
rect 465812 687012 465996 687176
rect 466212 687012 466370 687176
rect 468212 688212 468396 688376
rect 468612 688212 468796 688376
rect 468212 687812 468396 687976
rect 468612 687812 468796 687976
rect 468212 687412 468396 687576
rect 468612 687412 468796 687576
rect 468212 687012 468396 687176
rect 468622 687012 468806 687176
rect 415460 685408 415562 685516
rect 415820 685408 415922 685516
rect 415460 685168 415562 685276
rect 415820 685168 415922 685276
rect 467360 685404 467462 685512
rect 467720 685404 467822 685512
rect 467360 685164 467462 685272
rect 467720 685164 467822 685272
rect 66881 663007 66915 663109
rect 66986 663018 67068 663096
rect 74241 662809 74275 662911
rect 440260 657608 440362 657716
rect 440620 657608 440722 657716
rect 440260 657368 440362 657476
rect 440620 657368 440722 657476
rect 448860 657608 448962 657716
rect 449220 657608 449322 657716
rect 448860 657368 448962 657476
rect 449220 657368 449322 657476
rect 437812 656212 437996 656376
rect 438212 656212 438396 656376
rect 442412 656326 442596 656490
rect 442812 656326 442996 656490
rect 437812 655812 437996 655976
rect 438212 655812 438396 655976
rect 442412 655926 442596 656090
rect 442812 655926 442996 656090
rect 437812 655412 437996 655576
rect 438212 655412 438396 655576
rect 442412 655526 442596 655690
rect 442812 655526 442996 655690
rect 437812 655012 437996 655176
rect 438212 655012 438396 655176
rect 442412 655126 442596 655290
rect 442822 655126 443006 655290
rect 446212 656212 446396 656376
rect 446612 656212 446796 656376
rect 450812 656326 450996 656490
rect 451212 656326 451396 656490
rect 446212 655812 446396 655976
rect 446612 655812 446796 655976
rect 450814 655926 450996 656090
rect 451212 655926 451396 656090
rect 446212 655412 446396 655576
rect 446612 655412 446796 655576
rect 450814 655526 450996 655690
rect 451212 655526 451396 655690
rect 446212 655012 446396 655176
rect 446612 655012 446796 655176
rect 450814 655190 450996 655290
rect 450812 655126 450996 655190
rect 451222 655126 451406 655290
rect 440260 654608 440362 654716
rect 440620 654608 440722 654716
rect 440260 654368 440362 654476
rect 440620 654368 440722 654476
rect 448860 654608 448962 654716
rect 449220 654608 449322 654716
rect 448860 654368 448962 654476
rect 449220 654368 449322 654476
rect 134560 600104 134868 600344
rect 135160 600104 135468 600344
rect 135760 600104 136068 600344
rect 136360 600104 136668 600344
rect 136960 600104 137268 600344
rect 137560 600104 137868 600344
rect 138160 600104 138468 600344
rect 134006 599540 134086 599596
rect 134126 599540 134206 599596
rect 140406 599540 140486 599596
rect 140526 599540 140606 599596
rect 134006 599440 134086 599496
rect 134126 599440 134206 599496
rect 140406 599440 140486 599496
rect 140526 599440 140606 599496
rect 134398 598866 134592 599030
rect 134798 598866 134992 599030
rect 135198 598866 135392 599030
rect 135598 598866 135792 599030
rect 135998 598866 136192 599030
rect 136398 598866 136592 599030
rect 136798 598866 136992 599030
rect 137198 598866 137392 599030
rect 137598 598866 137792 599030
rect 137998 598866 138192 599030
rect 138398 598866 138592 599030
rect 138798 598866 138992 599030
rect 134398 598626 134592 598790
rect 134798 598626 134992 598790
rect 135198 598626 135392 598790
rect 135598 598626 135792 598790
rect 135998 598626 136192 598790
rect 136398 598626 136592 598790
rect 136798 598626 136992 598790
rect 137198 598626 137392 598790
rect 137598 598626 137792 598790
rect 137998 598626 138192 598790
rect 138398 598626 138592 598790
rect 138798 598626 138992 598790
rect 85560 586104 85868 586344
rect 86160 586104 86468 586344
rect 86760 586104 87068 586344
rect 87360 586104 87668 586344
rect 87960 586104 88268 586344
rect 88560 586104 88868 586344
rect 89160 586104 89468 586344
rect 424142 586174 424184 586416
rect 85006 585540 85086 585596
rect 85126 585540 85206 585596
rect 91406 585540 91486 585596
rect 91526 585540 91606 585596
rect 85006 585440 85086 585496
rect 85126 585440 85206 585496
rect 91406 585440 91486 585496
rect 91526 585440 91606 585496
rect 85398 584866 85592 585030
rect 85798 584866 85992 585030
rect 86198 584866 86392 585030
rect 86598 584866 86792 585030
rect 86998 584866 87192 585030
rect 87398 584866 87592 585030
rect 87798 584866 87992 585030
rect 88198 584866 88392 585030
rect 88598 584866 88792 585030
rect 88998 584866 89192 585030
rect 89398 584866 89592 585030
rect 89798 584866 89992 585030
rect 424132 584824 424174 585046
rect 85398 584626 85592 584790
rect 85798 584626 85992 584790
rect 86198 584626 86392 584790
rect 86598 584626 86792 584790
rect 86998 584626 87192 584790
rect 87398 584626 87592 584790
rect 87798 584626 87992 584790
rect 88198 584626 88392 584790
rect 88598 584626 88792 584790
rect 88998 584626 89192 584790
rect 89398 584626 89592 584790
rect 89798 584626 89992 584790
rect 101854 568504 102162 568744
rect 102454 568504 102762 568744
rect 103054 568504 103362 568744
rect 103654 568504 103962 568744
rect 104254 568504 104562 568744
rect 104854 568504 105162 568744
rect 105454 568504 105762 568744
rect 107560 568504 107868 568744
rect 108160 568504 108468 568744
rect 108760 568504 109068 568744
rect 109360 568504 109668 568744
rect 109960 568504 110268 568744
rect 110560 568504 110868 568744
rect 111160 568504 111468 568744
rect 102864 567740 102944 567796
rect 102984 567740 103064 567796
rect 104006 567740 104086 567796
rect 104126 567740 104206 567796
rect 102864 567640 102944 567696
rect 102984 567640 103064 567696
rect 104006 567640 104086 567696
rect 104126 567640 104206 567696
rect 107006 567740 107086 567796
rect 107126 567740 107206 567796
rect 113406 567788 113486 567844
rect 113526 567788 113606 567844
rect 107006 567640 107086 567696
rect 107126 567640 107206 567696
rect 113406 567688 113486 567744
rect 113526 567688 113606 567744
rect 101408 566904 101602 567068
rect 101808 566904 102002 567068
rect 102208 566904 102402 567068
rect 102608 566904 102802 567068
rect 103008 566904 103202 567068
rect 103408 566904 103602 567068
rect 103808 566904 104002 567068
rect 104208 566904 104402 567068
rect 104608 566904 104802 567068
rect 105008 566904 105202 567068
rect 105408 566904 105602 567068
rect 105808 566904 106002 567068
rect 101408 566664 101602 566828
rect 101808 566664 102002 566828
rect 102208 566664 102402 566828
rect 102608 566664 102802 566828
rect 103008 566664 103202 566828
rect 103408 566664 103602 566828
rect 103808 566664 104002 566828
rect 104208 566664 104402 566828
rect 104608 566664 104802 566828
rect 105008 566664 105202 566828
rect 105408 566664 105602 566828
rect 105808 566664 106002 566828
rect 107398 566866 107592 567030
rect 107798 567024 107908 567030
rect 107798 566866 107992 567024
rect 108198 566866 108392 567024
rect 108598 566866 108792 567024
rect 108998 566866 109192 567024
rect 109398 566866 109592 567024
rect 109798 566866 109992 567024
rect 110198 566866 110392 567030
rect 110598 566866 110792 567030
rect 110998 566866 111192 567030
rect 111398 566866 111592 567030
rect 111798 566866 111992 567030
rect 107398 566626 107592 566790
rect 107798 566626 107992 566790
rect 108198 566626 108392 566790
rect 108598 566626 108792 566790
rect 108998 566626 109192 566790
rect 109398 566626 109592 566790
rect 109798 566626 109992 566790
rect 110198 566626 110392 566790
rect 110598 566626 110792 566790
rect 110998 566626 111192 566790
rect 111398 566626 111592 566790
rect 111798 566626 111992 566790
<< metal1 >>
rect 116600 695294 118404 695994
rect 116600 694702 117144 695294
rect 117816 695206 118404 695294
rect 120132 695336 125206 695758
rect 117816 695109 118904 695206
rect 117816 695007 118843 695109
rect 118877 695007 118904 695109
rect 117816 694910 118904 695007
rect 118938 695164 119510 695166
rect 120132 695164 121002 695336
rect 118938 694978 121002 695164
rect 117816 694702 118404 694910
rect 116600 694138 118404 694702
rect 120132 694644 121002 694978
rect 121886 694644 123402 695336
rect 124286 694962 125206 695336
rect 126826 695396 128630 696096
rect 124286 694770 126154 694962
rect 126826 694940 127370 695396
rect 126190 694905 127370 694940
rect 126190 694803 126213 694905
rect 126247 694804 127370 694905
rect 128042 695308 128630 695396
rect 128042 695012 128634 695308
rect 128042 694804 128630 695012
rect 126247 694803 128630 694804
rect 126190 694792 128630 694803
rect 124286 694644 125206 694770
rect 120132 694286 125206 694644
rect 126826 694240 128630 694792
rect 467316 691416 467882 691454
rect 415416 691316 415982 691358
rect 415416 691208 415460 691316
rect 415562 691208 415820 691316
rect 415922 691208 415982 691316
rect 415416 691076 415982 691208
rect 415416 690968 415460 691076
rect 415562 690968 415820 691076
rect 415922 690968 415982 691076
rect 467316 691308 467360 691416
rect 467462 691308 467720 691416
rect 467822 691308 467882 691416
rect 467316 691176 467882 691308
rect 467316 691068 467360 691176
rect 467462 691068 467720 691176
rect 467822 691068 467882 691176
rect 467316 691026 467882 691068
rect 415416 690926 415982 690968
rect 413730 688376 414462 688608
rect 413730 688212 413812 688376
rect 413996 688212 414212 688376
rect 414396 688212 414462 688376
rect 413730 687976 414462 688212
rect 413730 687812 413812 687976
rect 413996 687812 414212 687976
rect 414396 687812 414462 687976
rect 413730 687576 414462 687812
rect 413730 687412 413812 687576
rect 413996 687412 414212 687576
rect 414396 687412 414462 687576
rect 413730 687176 414462 687412
rect 413730 687012 413812 687176
rect 413996 687012 414212 687176
rect 414396 687012 414462 687176
rect 413730 686944 414462 687012
rect 416130 688376 416866 688598
rect 416130 688212 416212 688376
rect 416396 688212 416612 688376
rect 416796 688212 416866 688376
rect 416130 687976 416866 688212
rect 416130 687812 416212 687976
rect 416396 687812 416612 687976
rect 416796 687812 416866 687976
rect 416130 687576 416866 687812
rect 416130 687412 416212 687576
rect 416396 687412 416612 687576
rect 416796 687412 416866 687576
rect 416130 687176 416866 687412
rect 416130 687012 416212 687176
rect 416396 687012 416622 687176
rect 416806 687012 416866 687176
rect 416130 686944 416866 687012
rect 465730 688376 466466 688608
rect 465730 688212 465812 688376
rect 465996 688212 466212 688376
rect 466396 688212 466466 688376
rect 465730 687976 466466 688212
rect 465730 687812 465812 687976
rect 465996 687812 466212 687976
rect 466396 687812 466466 687976
rect 465730 687576 466466 687812
rect 465730 687412 465812 687576
rect 465996 687412 466212 687576
rect 466396 687412 466466 687576
rect 465730 687176 466466 687412
rect 465730 687012 465812 687176
rect 465996 687012 466212 687176
rect 466396 687012 466466 687176
rect 465730 686944 466466 687012
rect 468130 688376 468866 688598
rect 468130 688212 468212 688376
rect 468396 688212 468612 688376
rect 468796 688212 468866 688376
rect 468130 687976 468866 688212
rect 468130 687812 468212 687976
rect 468396 687812 468612 687976
rect 468796 687812 468866 687976
rect 468130 687576 468866 687812
rect 468130 687412 468212 687576
rect 468396 687412 468612 687576
rect 468796 687412 468866 687576
rect 468130 687176 468866 687412
rect 468130 687012 468212 687176
rect 468396 687012 468622 687176
rect 468806 687012 468866 687176
rect 468130 686944 468866 687012
rect 415416 685516 415982 685558
rect 415416 685408 415460 685516
rect 415562 685408 415820 685516
rect 415922 685408 415982 685516
rect 415416 685276 415982 685408
rect 415416 685168 415460 685276
rect 415562 685168 415820 685276
rect 415922 685168 415982 685276
rect 415416 685126 415982 685168
rect 467316 685512 467882 685554
rect 467316 685404 467360 685512
rect 467462 685404 467720 685512
rect 467822 685404 467882 685512
rect 467316 685272 467882 685404
rect 467316 685164 467360 685272
rect 467462 685164 467720 685272
rect 467822 685164 467882 685272
rect 467316 685122 467882 685164
rect 64600 663294 66404 663994
rect 64600 662702 65144 663294
rect 65816 663206 66404 663294
rect 68132 663336 73206 663758
rect 65816 663109 66932 663206
rect 68132 663164 69002 663336
rect 65816 663007 66881 663109
rect 66915 663007 66932 663109
rect 65816 662910 66932 663007
rect 66976 663096 69002 663164
rect 66976 663018 66986 663096
rect 67068 663018 69002 663096
rect 66976 662978 69002 663018
rect 65816 662702 66404 662910
rect 64600 662138 66404 662702
rect 68132 662644 69002 662978
rect 69886 662644 71402 663336
rect 72286 662962 73206 663336
rect 74826 663396 76630 664096
rect 72286 662770 74184 662962
rect 74826 662940 75370 663396
rect 74220 662911 75370 662940
rect 74220 662809 74241 662911
rect 74275 662809 75370 662911
rect 74220 662804 75370 662809
rect 76042 663308 76630 663396
rect 76042 663012 76634 663308
rect 76042 662804 76630 663012
rect 74220 662792 76630 662804
rect 72286 662644 73206 662770
rect 68132 662286 73206 662644
rect 74826 662240 76630 662792
rect 440216 657716 440782 657758
rect 440216 657608 440260 657716
rect 440362 657608 440620 657716
rect 440722 657608 440782 657716
rect 440216 657476 440782 657608
rect 440216 657368 440260 657476
rect 440362 657368 440620 657476
rect 440722 657368 440782 657476
rect 440216 657328 440782 657368
rect 448816 657716 449382 657758
rect 448816 657608 448860 657716
rect 448962 657608 449220 657716
rect 449322 657608 449382 657716
rect 448816 657476 449382 657608
rect 448816 657368 448860 657476
rect 448962 657368 449220 657476
rect 449322 657368 449382 657476
rect 448816 657328 449382 657368
rect 437730 656376 438466 656608
rect 437730 656212 437812 656376
rect 437996 656212 438212 656376
rect 438396 656212 438466 656376
rect 437730 655976 438466 656212
rect 437730 655812 437812 655976
rect 437996 655812 438212 655976
rect 438396 655812 438466 655976
rect 437730 655576 438466 655812
rect 437730 655412 437812 655576
rect 437996 655412 438212 655576
rect 438396 655412 438466 655576
rect 437730 655176 438466 655412
rect 437730 655012 437812 655176
rect 437996 655012 438212 655176
rect 438396 655012 438466 655176
rect 442330 656490 443066 656712
rect 442330 656326 442412 656490
rect 442596 656326 442812 656490
rect 442996 656326 443066 656490
rect 442330 656090 443066 656326
rect 442330 655926 442412 656090
rect 442596 655926 442812 656090
rect 442996 655926 443066 656090
rect 442330 655690 443066 655926
rect 442330 655526 442412 655690
rect 442596 655526 442812 655690
rect 442996 655526 443066 655690
rect 442330 655290 443066 655526
rect 442330 655126 442412 655290
rect 442596 655126 442822 655290
rect 443006 655126 443066 655290
rect 442330 655058 443066 655126
rect 446130 656376 446866 656608
rect 446130 656212 446212 656376
rect 446396 656212 446612 656376
rect 446796 656212 446866 656376
rect 446130 655976 446866 656212
rect 446130 655812 446212 655976
rect 446396 655812 446612 655976
rect 446796 655812 446866 655976
rect 446130 655576 446866 655812
rect 446130 655412 446212 655576
rect 446396 655412 446612 655576
rect 446796 655412 446866 655576
rect 446130 655176 446866 655412
rect 437730 654944 438466 655012
rect 446130 655012 446212 655176
rect 446396 655012 446612 655176
rect 446796 655012 446866 655176
rect 450730 656490 451466 656712
rect 450730 656326 450812 656490
rect 450996 656326 451212 656490
rect 451396 656326 451466 656490
rect 450730 656090 451466 656326
rect 450730 655926 450812 656090
rect 450996 655926 451212 656090
rect 451396 655926 451466 656090
rect 450730 655690 451466 655926
rect 450730 655526 450812 655690
rect 450996 655526 451212 655690
rect 451396 655526 451466 655690
rect 450730 655290 451466 655526
rect 450730 655126 450812 655290
rect 450996 655126 451222 655290
rect 451406 655126 451466 655290
rect 450730 655058 451466 655126
rect 446130 654944 446866 655012
rect 440216 654716 440782 654758
rect 440216 654608 440260 654716
rect 440362 654608 440620 654716
rect 440722 654608 440782 654716
rect 440216 654476 440782 654608
rect 440216 654368 440260 654476
rect 440362 654368 440620 654476
rect 440722 654368 440782 654476
rect 440216 654328 440782 654368
rect 448816 654716 449382 654758
rect 448816 654608 448860 654716
rect 448962 654608 449220 654716
rect 449322 654608 449382 654716
rect 448816 654476 449382 654608
rect 448816 654368 448860 654476
rect 448962 654368 449220 654476
rect 449322 654368 449382 654476
rect 448816 654328 449382 654368
rect 134388 600344 139080 600454
rect 134388 600104 134560 600344
rect 134868 600104 135160 600344
rect 135468 600104 135760 600344
rect 136068 600104 136360 600344
rect 136668 600104 136960 600344
rect 137268 600104 137560 600344
rect 137868 600104 138160 600344
rect 138468 600104 139080 600344
rect 134388 600024 139080 600104
rect 134618 599942 135016 600024
rect 136144 599942 137882 600024
rect 134620 599830 135014 599942
rect 136150 599802 137878 599942
rect 133984 599596 134258 599606
rect 133984 599540 134006 599596
rect 134086 599540 134126 599596
rect 134206 599540 134258 599596
rect 133984 599496 134258 599540
rect 133984 599440 134006 599496
rect 134086 599440 134126 599496
rect 134206 599440 134258 599496
rect 133984 599410 134258 599440
rect 140384 599596 140628 599606
rect 140384 599540 140406 599596
rect 140486 599540 140526 599596
rect 140606 599540 140628 599596
rect 140384 599496 140628 599540
rect 140384 599440 140406 599496
rect 140486 599440 140526 599496
rect 140606 599440 140628 599496
rect 140384 599410 140628 599440
rect 134234 599060 134360 599078
rect 134602 599060 135002 599214
rect 136178 599060 138186 599252
rect 134234 599030 139092 599060
rect 134234 598866 134398 599030
rect 134592 598866 134798 599030
rect 134992 598866 135198 599030
rect 135392 598866 135598 599030
rect 135792 598866 135998 599030
rect 136192 598866 136398 599030
rect 136592 598866 136798 599030
rect 136992 598866 137198 599030
rect 137392 598866 137598 599030
rect 137792 598866 137998 599030
rect 138192 598866 138398 599030
rect 138592 598866 138798 599030
rect 138992 598866 139092 599030
rect 134234 598790 139092 598866
rect 134234 598626 134398 598790
rect 134592 598626 134798 598790
rect 134992 598626 135198 598790
rect 135392 598626 135598 598790
rect 135792 598626 135998 598790
rect 136192 598626 136398 598790
rect 136592 598626 136798 598790
rect 136992 598626 137198 598790
rect 137392 598626 137598 598790
rect 137792 598626 137998 598790
rect 138192 598626 138398 598790
rect 138592 598626 138798 598790
rect 138992 598626 139092 598790
rect 134234 598538 139092 598626
rect 134236 598260 139092 598538
rect 134234 597544 139096 598260
rect 134234 596998 134622 597544
rect 135400 596998 135822 597544
rect 136600 596998 137022 597544
rect 137800 596998 138222 597544
rect 139000 596998 139096 597544
rect 134234 596598 139096 596998
rect 416354 586782 417192 586912
rect 85388 586344 90080 586454
rect 85388 586104 85560 586344
rect 85868 586104 86160 586344
rect 86468 586104 86760 586344
rect 87068 586104 87360 586344
rect 87668 586104 87960 586344
rect 88268 586104 88560 586344
rect 88868 586104 89160 586344
rect 89468 586104 90080 586344
rect 416354 586394 416472 586782
rect 417092 586588 417192 586782
rect 417298 586588 417720 586590
rect 417092 586394 417970 586588
rect 425078 586450 428284 586452
rect 438104 586450 440896 586452
rect 441242 586450 441936 586452
rect 416354 586298 417970 586394
rect 416354 586296 417336 586298
rect 417712 586218 417970 586298
rect 424124 586446 428284 586450
rect 433144 586446 441936 586450
rect 424124 586416 441936 586446
rect 85388 586024 90080 586104
rect 85618 585788 86016 586024
rect 87144 585808 88882 586024
rect 417710 585916 418050 586218
rect 424124 586174 424142 586416
rect 424184 586394 441936 586416
rect 424184 586180 438974 586394
rect 441846 586214 441936 586394
rect 441846 586180 441958 586214
rect 424184 586174 441958 586180
rect 424124 586140 441958 586174
rect 425078 586138 441958 586140
rect 426680 586136 438282 586138
rect 426680 586132 433278 586136
rect 438896 586134 441958 586138
rect 426680 586126 428284 586132
rect 84984 585596 85258 585606
rect 84984 585540 85006 585596
rect 85086 585540 85126 585596
rect 85206 585540 85258 585596
rect 84984 585496 85258 585540
rect 84984 585440 85006 585496
rect 85086 585440 85126 585496
rect 85206 585440 85258 585496
rect 84984 585410 85258 585440
rect 91384 585596 91628 585606
rect 91384 585540 91406 585596
rect 91486 585540 91526 585596
rect 91606 585540 91628 585596
rect 91384 585496 91628 585540
rect 91384 585440 91406 585496
rect 91486 585440 91526 585496
rect 91606 585440 91628 585496
rect 91384 585410 91628 585440
rect 417624 585392 417840 585394
rect 85234 585076 85488 585078
rect 85632 585076 86000 585208
rect 87146 585076 88970 585218
rect 417066 585172 417284 585174
rect 416354 585170 417290 585172
rect 417624 585170 418062 585392
rect 416354 585098 418062 585170
rect 85234 585030 90092 585076
rect 85234 584866 85398 585030
rect 85592 584866 85798 585030
rect 85992 584866 86198 585030
rect 86392 584866 86598 585030
rect 86792 584866 86998 585030
rect 87192 584866 87398 585030
rect 87592 584866 87798 585030
rect 87992 584866 88198 585030
rect 88392 584866 88598 585030
rect 88792 584866 88998 585030
rect 89192 584866 89398 585030
rect 89592 584866 89798 585030
rect 89992 584866 90092 585030
rect 85234 584790 90092 584866
rect 85234 584626 85398 584790
rect 85592 584626 85798 584790
rect 85992 584626 86198 584790
rect 86392 584626 86598 584790
rect 86792 584626 86998 584790
rect 87192 584626 87398 584790
rect 87592 584626 87798 584790
rect 87992 584626 88198 584790
rect 88392 584626 88598 584790
rect 88792 584626 88998 584790
rect 89192 584626 89398 584790
rect 89592 584626 89798 584790
rect 89992 584626 90092 584790
rect 85234 584538 90092 584626
rect 416354 585072 417840 585098
rect 416354 584684 416472 585072
rect 417092 584876 417840 585072
rect 417092 584684 417186 584876
rect 417290 584874 417840 584876
rect 424118 585096 425178 585098
rect 426686 585096 450516 585098
rect 424118 585046 450516 585096
rect 417290 584872 417720 584874
rect 424118 584824 424132 585046
rect 424174 585042 450516 585046
rect 424174 584840 447368 585042
rect 450242 584840 450516 585042
rect 424174 584824 450516 584840
rect 424118 584792 450516 584824
rect 426686 584790 450516 584792
rect 416354 584586 417186 584684
rect 85236 584260 90092 584538
rect 85234 583544 90096 584260
rect 85234 582998 85622 583544
rect 86400 582998 86822 583544
rect 87600 582998 88022 583544
rect 88800 582998 89222 583544
rect 90000 582998 90096 583544
rect 85234 582598 90096 582998
rect 101682 568744 106034 568854
rect 101682 568504 101854 568744
rect 102162 568504 102454 568744
rect 102762 568504 103054 568744
rect 103362 568504 103654 568744
rect 103962 568504 104254 568744
rect 104562 568504 104854 568744
rect 105162 568504 105454 568744
rect 105762 568504 106034 568744
rect 101682 568424 106034 568504
rect 107388 568744 111740 568854
rect 107388 568504 107560 568744
rect 107868 568504 108160 568744
rect 108468 568504 108760 568744
rect 109068 568504 109360 568744
rect 109668 568504 109960 568744
rect 110268 568504 110560 568744
rect 110868 568504 111160 568744
rect 111468 568504 111740 568744
rect 107388 568424 111740 568504
rect 113384 567844 113620 567854
rect 102842 567796 103076 567806
rect 102842 567740 102864 567796
rect 102944 567740 102984 567796
rect 103064 567740 103076 567796
rect 102842 567696 103076 567740
rect 102842 567640 102864 567696
rect 102944 567640 102984 567696
rect 103064 567640 103076 567696
rect 102842 567610 103076 567640
rect 103986 567796 104220 567806
rect 103986 567740 104006 567796
rect 104086 567740 104126 567796
rect 104206 567740 104220 567796
rect 103986 567696 104220 567740
rect 103986 567640 104006 567696
rect 104086 567640 104126 567696
rect 104206 567640 104220 567696
rect 103986 567610 104220 567640
rect 106984 567796 107220 567806
rect 106984 567740 107006 567796
rect 107086 567740 107126 567796
rect 107206 567740 107220 567796
rect 106984 567696 107220 567740
rect 106984 567640 107006 567696
rect 107086 567640 107126 567696
rect 107206 567640 107220 567696
rect 113384 567788 113406 567844
rect 113486 567788 113526 567844
rect 113606 567788 113620 567844
rect 113384 567744 113620 567788
rect 113384 567688 113406 567744
rect 113486 567688 113526 567744
rect 113606 567688 113620 567744
rect 113384 567658 113620 567688
rect 106984 567610 107220 567640
rect 101244 567114 101498 567116
rect 102880 567114 103904 567454
rect 101244 567068 106102 567114
rect 101244 566904 101408 567068
rect 101602 566904 101808 567068
rect 102002 566904 102208 567068
rect 102402 566904 102608 567068
rect 102802 566904 103008 567068
rect 103202 566904 103408 567068
rect 103602 566904 103808 567068
rect 104002 566904 104208 567068
rect 104402 566904 104608 567068
rect 104802 566904 105008 567068
rect 105202 566904 105408 567068
rect 105602 566904 105808 567068
rect 106002 566904 106102 567068
rect 101244 566828 106102 566904
rect 101244 566664 101408 566828
rect 101602 566664 101808 566828
rect 102002 566664 102208 566828
rect 102402 566664 102608 566828
rect 102802 566664 103008 566828
rect 103202 566664 103408 566828
rect 103602 566664 103808 566828
rect 104002 566664 104208 566828
rect 104402 566664 104608 566828
rect 104802 566664 105008 566828
rect 105202 566664 105408 566828
rect 105602 566664 105808 566828
rect 106002 566664 106102 566828
rect 101244 566576 106102 566664
rect 101246 566298 106102 566576
rect 107234 567076 107488 567078
rect 107234 567030 112092 567076
rect 107234 566866 107398 567030
rect 107592 566866 107798 567030
rect 107908 567024 110198 567030
rect 107992 566866 108198 567024
rect 108392 566866 108598 567024
rect 108792 566866 108998 567024
rect 109192 566866 109398 567024
rect 109592 566866 109798 567024
rect 109992 566866 110198 567024
rect 110392 566866 110598 567030
rect 110792 566866 110998 567030
rect 111192 566866 111398 567030
rect 111592 566866 111798 567030
rect 111992 566866 112092 567030
rect 107234 566790 112092 566866
rect 107234 566626 107398 566790
rect 107592 566626 107798 566790
rect 107992 566626 108198 566790
rect 108392 566626 108598 566790
rect 108792 566626 108998 566790
rect 109192 566626 109398 566790
rect 109592 566626 109798 566790
rect 109992 566626 110198 566790
rect 110392 566626 110598 566790
rect 110792 566626 110998 566790
rect 111192 566626 111398 566790
rect 111592 566626 111798 566790
rect 111992 566626 112092 566790
rect 107234 566538 112092 566626
rect 101244 565582 106106 566298
rect 107236 566260 112092 566538
rect 101244 565036 101632 565582
rect 102410 565036 102832 565582
rect 103610 565036 104032 565582
rect 104810 565036 105232 565582
rect 106010 565036 106106 565582
rect 101244 564636 106106 565036
rect 107234 565544 112096 566260
rect 107234 564998 107622 565544
rect 108400 564998 108822 565544
rect 109600 564998 110022 565544
rect 110800 564998 111222 565544
rect 112000 564998 112096 565544
rect 107234 564598 112096 564998
<< via1 >>
rect 117144 694702 117816 695294
rect 121002 694644 121886 695336
rect 123402 694644 124286 695336
rect 127370 694804 128042 695396
rect 415460 691208 415562 691316
rect 415820 691208 415922 691316
rect 415460 690968 415562 691076
rect 415820 690968 415922 691076
rect 467360 691308 467462 691416
rect 467720 691308 467822 691416
rect 467360 691068 467462 691176
rect 467720 691068 467822 691176
rect 413812 688212 413996 688376
rect 414212 688212 414394 688376
rect 414394 688212 414396 688376
rect 413812 687812 413996 687976
rect 414212 687812 414394 687976
rect 414394 687812 414396 687976
rect 413812 687412 413996 687576
rect 414212 687412 414394 687576
rect 414394 687412 414396 687576
rect 413812 687012 413996 687176
rect 414212 687012 414394 687176
rect 414394 687012 414396 687176
rect 416212 688212 416396 688376
rect 416612 688212 416796 688376
rect 416212 687812 416396 687976
rect 416612 687812 416796 687976
rect 416212 687412 416396 687576
rect 416612 687412 416796 687576
rect 416212 687012 416396 687176
rect 416622 687012 416806 687176
rect 465812 688212 465996 688376
rect 466212 688212 466370 688376
rect 466370 688212 466396 688376
rect 465812 687812 465996 687976
rect 466212 687812 466370 687976
rect 466370 687812 466396 687976
rect 465812 687412 465996 687576
rect 466212 687412 466370 687576
rect 466370 687412 466396 687576
rect 465812 687012 465996 687176
rect 466212 687012 466370 687176
rect 466370 687012 466396 687176
rect 468212 688212 468396 688376
rect 468612 688212 468796 688376
rect 468212 687812 468396 687976
rect 468612 687812 468796 687976
rect 468212 687412 468396 687576
rect 468612 687412 468796 687576
rect 468212 687012 468396 687176
rect 468622 687012 468806 687176
rect 415460 685408 415562 685516
rect 415820 685408 415922 685516
rect 415460 685168 415562 685276
rect 415820 685168 415922 685276
rect 467360 685404 467462 685512
rect 467720 685404 467822 685512
rect 467360 685164 467462 685272
rect 467720 685164 467822 685272
rect 65144 662702 65816 663294
rect 69002 662644 69886 663336
rect 71402 662644 72286 663336
rect 75370 662804 76042 663396
rect 440260 657608 440362 657716
rect 440620 657608 440722 657716
rect 440260 657368 440362 657476
rect 440620 657368 440722 657476
rect 448860 657608 448962 657716
rect 449220 657608 449322 657716
rect 448860 657368 448962 657476
rect 449220 657368 449322 657476
rect 437812 656212 437996 656376
rect 438212 656212 438396 656376
rect 437812 655812 437996 655976
rect 438212 655812 438396 655976
rect 437812 655412 437996 655576
rect 438212 655412 438396 655576
rect 437812 655012 437996 655176
rect 438212 655012 438396 655176
rect 442412 656326 442596 656490
rect 442812 656326 442996 656490
rect 442412 655926 442596 656090
rect 442812 655926 442996 656090
rect 442412 655526 442596 655690
rect 442812 655526 442996 655690
rect 442412 655126 442596 655290
rect 442822 655126 443006 655290
rect 446212 656212 446396 656376
rect 446612 656212 446796 656376
rect 446212 655812 446396 655976
rect 446612 655812 446796 655976
rect 446212 655412 446396 655576
rect 446612 655412 446796 655576
rect 446212 655012 446396 655176
rect 446612 655012 446796 655176
rect 450812 656326 450996 656490
rect 451212 656326 451396 656490
rect 450812 655926 450814 656090
rect 450814 655926 450996 656090
rect 451212 655926 451396 656090
rect 450812 655526 450814 655690
rect 450814 655526 450996 655690
rect 451212 655526 451396 655690
rect 450812 655190 450814 655290
rect 450814 655190 450996 655290
rect 450812 655126 450996 655190
rect 451222 655126 451406 655290
rect 440260 654608 440362 654716
rect 440620 654608 440722 654716
rect 440260 654368 440362 654476
rect 440620 654368 440722 654476
rect 448860 654608 448962 654716
rect 449220 654608 449322 654716
rect 448860 654368 448962 654476
rect 449220 654368 449322 654476
rect 134560 600104 134868 600344
rect 135160 600104 135468 600344
rect 135760 600104 136068 600344
rect 136360 600104 136668 600344
rect 136960 600104 137268 600344
rect 137560 600104 137868 600344
rect 138160 600104 138468 600344
rect 134006 599540 134086 599596
rect 134126 599540 134206 599596
rect 134006 599440 134086 599496
rect 134126 599440 134206 599496
rect 140406 599540 140486 599596
rect 140526 599540 140606 599596
rect 140406 599440 140486 599496
rect 140526 599440 140606 599496
rect 134622 596998 135400 597544
rect 135822 596998 136600 597544
rect 137022 596998 137800 597544
rect 138222 596998 139000 597544
rect 85560 586104 85868 586344
rect 86160 586104 86468 586344
rect 86760 586104 87068 586344
rect 87360 586104 87668 586344
rect 87960 586104 88268 586344
rect 88560 586104 88868 586344
rect 89160 586104 89468 586344
rect 416472 586394 417092 586782
rect 438974 586180 441846 586394
rect 85006 585540 85086 585596
rect 85126 585540 85206 585596
rect 85006 585440 85086 585496
rect 85126 585440 85206 585496
rect 91406 585540 91486 585596
rect 91526 585540 91606 585596
rect 91406 585440 91486 585496
rect 91526 585440 91606 585496
rect 416472 584684 417092 585072
rect 447368 584840 450242 585042
rect 85622 582998 86400 583544
rect 86822 582998 87600 583544
rect 88022 582998 88800 583544
rect 89222 582998 90000 583544
rect 101854 568504 102162 568744
rect 102454 568504 102762 568744
rect 103054 568504 103362 568744
rect 103654 568504 103962 568744
rect 104254 568504 104562 568744
rect 104854 568504 105162 568744
rect 105454 568504 105762 568744
rect 107560 568504 107868 568744
rect 108160 568504 108468 568744
rect 108760 568504 109068 568744
rect 109360 568504 109668 568744
rect 109960 568504 110268 568744
rect 110560 568504 110868 568744
rect 111160 568504 111468 568744
rect 102864 567740 102944 567796
rect 102984 567740 103064 567796
rect 102864 567640 102944 567696
rect 102984 567640 103064 567696
rect 104006 567740 104086 567796
rect 104126 567740 104206 567796
rect 104006 567640 104086 567696
rect 104126 567640 104206 567696
rect 107006 567740 107086 567796
rect 107126 567740 107206 567796
rect 107006 567640 107086 567696
rect 107126 567640 107206 567696
rect 113406 567788 113486 567844
rect 113526 567788 113606 567844
rect 113406 567688 113486 567744
rect 113526 567688 113606 567744
rect 101632 565036 102410 565582
rect 102832 565036 103610 565582
rect 104032 565036 104810 565582
rect 105232 565036 106010 565582
rect 107622 564998 108400 565544
rect 108822 564998 109600 565544
rect 110022 564998 110800 565544
rect 111222 564998 112000 565544
<< metal2 >>
rect 116600 695398 118404 695994
rect 116600 694620 117052 695398
rect 117904 694620 118404 695398
rect 116600 694138 118404 694620
rect 120132 695502 125206 695758
rect 120132 694490 120888 695502
rect 122028 694490 123288 695502
rect 124428 694490 125206 695502
rect 120132 694286 125206 694490
rect 126826 695500 128630 696096
rect 126826 694722 127278 695500
rect 128130 694722 128630 695500
rect 126826 694240 128630 694722
rect 467316 691416 467882 691454
rect 415416 691316 415982 691358
rect 415416 691208 415460 691316
rect 415562 691208 415820 691316
rect 415922 691208 415982 691316
rect 415416 691076 415982 691208
rect 415416 690968 415460 691076
rect 415562 690968 415820 691076
rect 415922 690968 415982 691076
rect 467316 691308 467360 691416
rect 467462 691308 467720 691416
rect 467822 691308 467882 691416
rect 467316 691176 467882 691308
rect 467316 691068 467360 691176
rect 467462 691068 467720 691176
rect 467822 691068 467882 691176
rect 467316 691026 467882 691068
rect 415416 690926 415982 690968
rect 413730 688376 414462 688608
rect 413730 688212 413812 688376
rect 413996 688212 414212 688376
rect 414396 688212 414462 688376
rect 413730 687976 414462 688212
rect 413730 687812 413812 687976
rect 413996 687812 414212 687976
rect 414396 687812 414462 687976
rect 413730 687576 414462 687812
rect 413730 687412 413812 687576
rect 413996 687412 414212 687576
rect 414396 687412 414462 687576
rect 413730 687176 414462 687412
rect 413730 687012 413812 687176
rect 413996 687012 414212 687176
rect 414396 687012 414462 687176
rect 413730 686944 414462 687012
rect 416130 688376 416866 688598
rect 416130 688212 416212 688376
rect 416396 688212 416612 688376
rect 416796 688212 416866 688376
rect 416130 687976 416866 688212
rect 416130 687812 416212 687976
rect 416396 687812 416612 687976
rect 416796 687812 416866 687976
rect 416130 687576 416866 687812
rect 416130 687412 416212 687576
rect 416396 687412 416612 687576
rect 416796 687412 416866 687576
rect 416130 687176 416866 687412
rect 416130 687012 416212 687176
rect 416396 687012 416622 687176
rect 416806 687012 416866 687176
rect 416130 686944 416866 687012
rect 465730 688376 466466 688608
rect 465730 688212 465812 688376
rect 465996 688212 466212 688376
rect 466396 688212 466466 688376
rect 465730 687976 466466 688212
rect 465730 687812 465812 687976
rect 465996 687812 466212 687976
rect 466396 687812 466466 687976
rect 465730 687576 466466 687812
rect 465730 687412 465812 687576
rect 465996 687412 466212 687576
rect 466396 687412 466466 687576
rect 465730 687176 466466 687412
rect 465730 687012 465812 687176
rect 465996 687012 466212 687176
rect 466396 687012 466466 687176
rect 465730 686944 466466 687012
rect 468130 688376 468866 688598
rect 468130 688212 468212 688376
rect 468396 688212 468612 688376
rect 468796 688212 468866 688376
rect 468130 687976 468866 688212
rect 468130 687812 468212 687976
rect 468396 687812 468612 687976
rect 468796 687812 468866 687976
rect 468130 687576 468866 687812
rect 468130 687412 468212 687576
rect 468396 687412 468612 687576
rect 468796 687412 468866 687576
rect 468130 687176 468866 687412
rect 468130 687012 468212 687176
rect 468396 687012 468622 687176
rect 468806 687012 468866 687176
rect 468130 686944 468866 687012
rect 415416 685516 415982 685558
rect 415416 685408 415460 685516
rect 415562 685408 415820 685516
rect 415922 685408 415982 685516
rect 415416 685276 415982 685408
rect 415416 685168 415460 685276
rect 415562 685168 415820 685276
rect 415922 685168 415982 685276
rect 415416 685126 415982 685168
rect 467316 685512 467882 685554
rect 467316 685404 467360 685512
rect 467462 685404 467720 685512
rect 467822 685404 467882 685512
rect 467316 685272 467882 685404
rect 467316 685164 467360 685272
rect 467462 685164 467720 685272
rect 467822 685164 467882 685272
rect 467316 685122 467882 685164
rect 64600 663398 66404 663994
rect 64600 662620 65052 663398
rect 65904 662620 66404 663398
rect 64600 662138 66404 662620
rect 68132 663502 73206 663758
rect 68132 662490 68888 663502
rect 70028 662490 71288 663502
rect 72428 662490 73206 663502
rect 68132 662286 73206 662490
rect 74826 663500 76630 664096
rect 74826 662722 75278 663500
rect 76130 662722 76630 663500
rect 74826 662240 76630 662722
rect 440216 657716 440782 657758
rect 440216 657608 440260 657716
rect 440362 657608 440620 657716
rect 440722 657608 440782 657716
rect 440216 657476 440782 657608
rect 440216 657368 440260 657476
rect 440362 657368 440620 657476
rect 440722 657368 440782 657476
rect 440216 657328 440782 657368
rect 448816 657716 449382 657758
rect 448816 657608 448860 657716
rect 448962 657608 449220 657716
rect 449322 657608 449382 657716
rect 448816 657476 449382 657608
rect 448816 657368 448860 657476
rect 448962 657368 449220 657476
rect 449322 657368 449382 657476
rect 448816 657328 449382 657368
rect 437730 656376 438466 656608
rect 437730 656212 437812 656376
rect 437996 656212 438212 656376
rect 438396 656212 438466 656376
rect 437730 655976 438466 656212
rect 437730 655812 437812 655976
rect 437996 655812 438212 655976
rect 438396 655812 438466 655976
rect 437730 655576 438466 655812
rect 437730 655412 437812 655576
rect 437996 655412 438212 655576
rect 438396 655412 438466 655576
rect 437730 655176 438466 655412
rect 437730 655012 437812 655176
rect 437996 655012 438212 655176
rect 438396 655012 438466 655176
rect 442330 656490 443066 656712
rect 442330 656326 442412 656490
rect 442596 656326 442812 656490
rect 442996 656326 443066 656490
rect 442330 656090 443066 656326
rect 442330 655926 442412 656090
rect 442596 655926 442812 656090
rect 442996 655926 443066 656090
rect 442330 655690 443066 655926
rect 442330 655526 442412 655690
rect 442596 655526 442812 655690
rect 442996 655526 443066 655690
rect 442330 655290 443066 655526
rect 442330 655126 442412 655290
rect 442596 655126 442822 655290
rect 443006 655126 443066 655290
rect 442330 655058 443066 655126
rect 446130 656376 446866 656608
rect 446130 656212 446212 656376
rect 446396 656212 446612 656376
rect 446796 656212 446866 656376
rect 446130 655976 446866 656212
rect 446130 655812 446212 655976
rect 446396 655812 446612 655976
rect 446796 655812 446866 655976
rect 446130 655576 446866 655812
rect 446130 655412 446212 655576
rect 446396 655412 446612 655576
rect 446796 655412 446866 655576
rect 446130 655176 446866 655412
rect 437730 654944 438466 655012
rect 446130 655012 446212 655176
rect 446396 655012 446612 655176
rect 446796 655012 446866 655176
rect 450730 656490 451466 656712
rect 450730 656326 450812 656490
rect 450996 656326 451212 656490
rect 451396 656326 451466 656490
rect 450730 656090 451466 656326
rect 450730 655926 450812 656090
rect 450996 655926 451212 656090
rect 451396 655926 451466 656090
rect 450730 655690 451466 655926
rect 450730 655526 450812 655690
rect 450996 655526 451212 655690
rect 451396 655526 451466 655690
rect 450730 655290 451466 655526
rect 450730 655126 450812 655290
rect 450996 655126 451222 655290
rect 451406 655126 451466 655290
rect 450730 655058 451466 655126
rect 446130 654944 446866 655012
rect 440216 654716 440782 654758
rect 440216 654608 440260 654716
rect 440362 654608 440620 654716
rect 440722 654608 440782 654716
rect 440216 654476 440782 654608
rect 440216 654368 440260 654476
rect 440362 654368 440620 654476
rect 440722 654368 440782 654476
rect 440216 654328 440782 654368
rect 448816 654716 449382 654758
rect 448816 654608 448860 654716
rect 448962 654608 449220 654716
rect 449322 654608 449382 654716
rect 448816 654476 449382 654608
rect 448816 654368 448860 654476
rect 448962 654368 449220 654476
rect 449322 654368 449382 654476
rect 448816 654328 449382 654368
rect 134388 600344 139080 600454
rect 134388 600104 134560 600344
rect 134868 600104 135160 600344
rect 135468 600104 135760 600344
rect 136068 600104 136360 600344
rect 136668 600104 136960 600344
rect 137268 600104 137560 600344
rect 137868 600104 138160 600344
rect 138468 600104 139080 600344
rect 134388 600024 139080 600104
rect 133984 599596 134258 599606
rect 133984 599540 134006 599596
rect 134086 599540 134126 599596
rect 134206 599540 134258 599596
rect 133984 599496 134258 599540
rect 133984 599440 134006 599496
rect 134086 599440 134126 599496
rect 134206 599440 134258 599496
rect 133984 599410 134258 599440
rect 140384 599596 140628 599606
rect 140384 599540 140406 599596
rect 140486 599540 140526 599596
rect 140606 599540 140628 599596
rect 140384 599496 140628 599540
rect 140384 599440 140406 599496
rect 140486 599440 140526 599496
rect 140606 599440 140628 599496
rect 140384 599410 140628 599440
rect 134234 597544 139146 597958
rect 134234 596998 134622 597544
rect 135400 596998 135822 597544
rect 136600 596998 137022 597544
rect 137800 596998 138222 597544
rect 139000 596998 139146 597544
rect 134234 596602 139146 596998
rect 416354 586782 417192 586912
rect 85388 586344 90080 586454
rect 85388 586104 85560 586344
rect 85868 586104 86160 586344
rect 86468 586104 86760 586344
rect 87068 586104 87360 586344
rect 87668 586104 87960 586344
rect 88268 586104 88560 586344
rect 88868 586104 89160 586344
rect 89468 586104 90080 586344
rect 416354 586394 416472 586782
rect 417092 586394 417192 586782
rect 416354 586296 417192 586394
rect 438926 586394 441902 586434
rect 438926 586180 438974 586394
rect 441846 586180 441902 586394
rect 438926 586136 441902 586180
rect 85388 586024 90080 586104
rect 415786 585612 416282 585710
rect 415786 585608 417420 585612
rect 84984 585596 85258 585606
rect 84984 585540 85006 585596
rect 85086 585540 85126 585596
rect 85206 585540 85258 585596
rect 84984 585496 85258 585540
rect 84984 585440 85006 585496
rect 85086 585440 85126 585496
rect 85206 585440 85258 585496
rect 84984 585410 85258 585440
rect 91384 585596 91628 585606
rect 91384 585540 91406 585596
rect 91486 585540 91526 585596
rect 91606 585540 91628 585596
rect 91384 585496 91628 585540
rect 91384 585440 91406 585496
rect 91486 585440 91526 585496
rect 91606 585440 91628 585496
rect 91384 585410 91628 585440
rect 415786 585422 415878 585608
rect 416190 585422 417420 585608
rect 415786 585412 417420 585422
rect 415786 585344 416282 585412
rect 416354 585072 417186 585172
rect 416354 584684 416472 585072
rect 417092 584684 417186 585072
rect 447352 585042 450258 585064
rect 447352 584840 447368 585042
rect 450242 584840 450258 585042
rect 447352 584820 450258 584840
rect 416354 584586 417186 584684
rect 85234 583544 90146 583958
rect 85234 582998 85622 583544
rect 86400 582998 86822 583544
rect 87600 582998 88022 583544
rect 88800 582998 89222 583544
rect 90000 582998 90146 583544
rect 85234 582602 90146 582998
rect 101682 568744 106034 568854
rect 101682 568504 101854 568744
rect 102162 568504 102454 568744
rect 102762 568504 103054 568744
rect 103362 568504 103654 568744
rect 103962 568504 104254 568744
rect 104562 568504 104854 568744
rect 105162 568504 105454 568744
rect 105762 568504 106034 568744
rect 101682 568424 106034 568504
rect 107388 568744 111740 568854
rect 107388 568504 107560 568744
rect 107868 568504 108160 568744
rect 108468 568504 108760 568744
rect 109068 568504 109360 568744
rect 109668 568504 109960 568744
rect 110268 568504 110560 568744
rect 110868 568504 111160 568744
rect 111468 568504 111740 568744
rect 107388 568424 111740 568504
rect 113384 567844 113620 567854
rect 102842 567796 103076 567806
rect 102842 567740 102864 567796
rect 102944 567740 102984 567796
rect 103064 567740 103076 567796
rect 102842 567696 103076 567740
rect 102842 567640 102864 567696
rect 102944 567640 102984 567696
rect 103064 567640 103076 567696
rect 102842 567610 103076 567640
rect 103986 567796 104220 567806
rect 103986 567740 104006 567796
rect 104086 567740 104126 567796
rect 104206 567740 104220 567796
rect 103986 567696 104220 567740
rect 103986 567640 104006 567696
rect 104086 567640 104126 567696
rect 104206 567640 104220 567696
rect 103986 567610 104220 567640
rect 106984 567796 107220 567806
rect 106984 567740 107006 567796
rect 107086 567740 107126 567796
rect 107206 567740 107220 567796
rect 106984 567696 107220 567740
rect 106984 567640 107006 567696
rect 107086 567640 107126 567696
rect 107206 567640 107220 567696
rect 113384 567788 113406 567844
rect 113486 567788 113526 567844
rect 113606 567788 113620 567844
rect 113384 567744 113620 567788
rect 113384 567688 113406 567744
rect 113486 567688 113526 567744
rect 113606 567688 113620 567744
rect 113384 567658 113620 567688
rect 106984 567610 107220 567640
rect 101244 565582 106156 565996
rect 101244 565036 101632 565582
rect 102410 565036 102832 565582
rect 103610 565036 104032 565582
rect 104810 565036 105232 565582
rect 106010 565036 106156 565582
rect 101244 564640 106156 565036
rect 107234 565544 112146 565958
rect 107234 564998 107622 565544
rect 108400 564998 108822 565544
rect 109600 564998 110022 565544
rect 110800 564998 111222 565544
rect 112000 564998 112146 565544
rect 107234 564602 112146 564998
rect 524 -800 636 480
rect 1706 -800 1818 480
rect 2888 -800 3000 480
rect 4070 -800 4182 480
rect 5252 -800 5364 480
rect 6434 -800 6546 480
rect 7616 -800 7728 480
rect 8798 -800 8910 480
rect 9980 -800 10092 480
rect 11162 -800 11274 480
rect 12344 -800 12456 480
rect 13526 -800 13638 480
rect 14708 -800 14820 480
rect 15890 -800 16002 480
rect 17072 -800 17184 480
rect 18254 -800 18366 480
rect 19436 -800 19548 480
rect 20618 -800 20730 480
rect 21800 -800 21912 480
rect 22982 -800 23094 480
rect 24164 -800 24276 480
rect 25346 -800 25458 480
rect 26528 -800 26640 480
rect 27710 -800 27822 480
rect 28892 -800 29004 480
rect 30074 -800 30186 480
rect 31256 -800 31368 480
rect 32438 -800 32550 480
rect 33620 -800 33732 480
rect 34802 -800 34914 480
rect 35984 -800 36096 480
rect 37166 -800 37278 480
rect 38348 -800 38460 480
rect 39530 -800 39642 480
rect 40712 -800 40824 480
rect 41894 -800 42006 480
rect 43076 -800 43188 480
rect 44258 -800 44370 480
rect 45440 -800 45552 480
rect 46622 -800 46734 480
rect 47804 -800 47916 480
rect 48986 -800 49098 480
rect 50168 -800 50280 480
rect 51350 -800 51462 480
rect 52532 -800 52644 480
rect 53714 -800 53826 480
rect 54896 -800 55008 480
rect 56078 -800 56190 480
rect 57260 -800 57372 480
rect 58442 -800 58554 480
rect 59624 -800 59736 480
rect 60806 -800 60918 480
rect 61988 -800 62100 480
rect 63170 -800 63282 480
rect 64352 -800 64464 480
rect 65534 -800 65646 480
rect 66716 -800 66828 480
rect 67898 -800 68010 480
rect 69080 -800 69192 480
rect 70262 -800 70374 480
rect 71444 -800 71556 480
rect 72626 -800 72738 480
rect 73808 -800 73920 480
rect 74990 -800 75102 480
rect 76172 -800 76284 480
rect 77354 -800 77466 480
rect 78536 -800 78648 480
rect 79718 -800 79830 480
rect 80900 -800 81012 480
rect 82082 -800 82194 480
rect 83264 -800 83376 480
rect 84446 -800 84558 480
rect 85628 -800 85740 480
rect 86810 -800 86922 480
rect 87992 -800 88104 480
rect 89174 -800 89286 480
rect 90356 -800 90468 480
rect 91538 -800 91650 480
rect 92720 -800 92832 480
rect 93902 -800 94014 480
rect 95084 -800 95196 480
rect 96266 -800 96378 480
rect 97448 -800 97560 480
rect 98630 -800 98742 480
rect 99812 -800 99924 480
rect 100994 -800 101106 480
rect 102176 -800 102288 480
rect 103358 -800 103470 480
rect 104540 -800 104652 480
rect 105722 -800 105834 480
rect 106904 -800 107016 480
rect 108086 -800 108198 480
rect 109268 -800 109380 480
rect 110450 -800 110562 480
rect 111632 -800 111744 480
rect 112814 -800 112926 480
rect 113996 -800 114108 480
rect 115178 -800 115290 480
rect 116360 -800 116472 480
rect 117542 -800 117654 480
rect 118724 -800 118836 480
rect 119906 -800 120018 480
rect 121088 -800 121200 480
rect 122270 -800 122382 480
rect 123452 -800 123564 480
rect 124634 -800 124746 480
rect 125816 -800 125928 480
rect 126998 -800 127110 480
rect 128180 -800 128292 480
rect 129362 -800 129474 480
rect 130544 -800 130656 480
rect 131726 -800 131838 480
rect 132908 -800 133020 480
rect 134090 -800 134202 480
rect 135272 -800 135384 480
rect 136454 -800 136566 480
rect 137636 -800 137748 480
rect 138818 -800 138930 480
rect 140000 -800 140112 480
rect 141182 -800 141294 480
rect 142364 -800 142476 480
rect 143546 -800 143658 480
rect 144728 -800 144840 480
rect 145910 -800 146022 480
rect 147092 -800 147204 480
rect 148274 -800 148386 480
rect 149456 -800 149568 480
rect 150638 -800 150750 480
rect 151820 -800 151932 480
rect 153002 -800 153114 480
rect 154184 -800 154296 480
rect 155366 -800 155478 480
rect 156548 -800 156660 480
rect 157730 -800 157842 480
rect 158912 -800 159024 480
rect 160094 -800 160206 480
rect 161276 -800 161388 480
rect 162458 -800 162570 480
rect 163640 -800 163752 480
rect 164822 -800 164934 480
rect 166004 -800 166116 480
rect 167186 -800 167298 480
rect 168368 -800 168480 480
rect 169550 -800 169662 480
rect 170732 -800 170844 480
rect 171914 -800 172026 480
rect 173096 -800 173208 480
rect 174278 -800 174390 480
rect 175460 -800 175572 480
rect 176642 -800 176754 480
rect 177824 -800 177936 480
rect 179006 -800 179118 480
rect 180188 -800 180300 480
rect 181370 -800 181482 480
rect 182552 -800 182664 480
rect 183734 -800 183846 480
rect 184916 -800 185028 480
rect 186098 -800 186210 480
rect 187280 -800 187392 480
rect 188462 -800 188574 480
rect 189644 -800 189756 480
rect 190826 -800 190938 480
rect 192008 -800 192120 480
rect 193190 -800 193302 480
rect 194372 -800 194484 480
rect 195554 -800 195666 480
rect 196736 -800 196848 480
rect 197918 -800 198030 480
rect 199100 -800 199212 480
rect 200282 -800 200394 480
rect 201464 -800 201576 480
rect 202646 -800 202758 480
rect 203828 -800 203940 480
rect 205010 -800 205122 480
rect 206192 -800 206304 480
rect 207374 -800 207486 480
rect 208556 -800 208668 480
rect 209738 -800 209850 480
rect 210920 -800 211032 480
rect 212102 -800 212214 480
rect 213284 -800 213396 480
rect 214466 -800 214578 480
rect 215648 -800 215760 480
rect 216830 -800 216942 480
rect 218012 -800 218124 480
rect 219194 -800 219306 480
rect 220376 -800 220488 480
rect 221558 -800 221670 480
rect 222740 -800 222852 480
rect 223922 -800 224034 480
rect 225104 -800 225216 480
rect 226286 -800 226398 480
rect 227468 -800 227580 480
rect 228650 -800 228762 480
rect 229832 -800 229944 480
rect 231014 -800 231126 480
rect 232196 -800 232308 480
rect 233378 -800 233490 480
rect 234560 -800 234672 480
rect 235742 -800 235854 480
rect 236924 -800 237036 480
rect 238106 -800 238218 480
rect 239288 -800 239400 480
rect 240470 -800 240582 480
rect 241652 -800 241764 480
rect 242834 -800 242946 480
rect 244016 -800 244128 480
rect 245198 -800 245310 480
rect 246380 -800 246492 480
rect 247562 -800 247674 480
rect 248744 -800 248856 480
rect 249926 -800 250038 480
rect 251108 -800 251220 480
rect 252290 -800 252402 480
rect 253472 -800 253584 480
rect 254654 -800 254766 480
rect 255836 -800 255948 480
rect 257018 -800 257130 480
rect 258200 -800 258312 480
rect 259382 -800 259494 480
rect 260564 -800 260676 480
rect 261746 -800 261858 480
rect 262928 -800 263040 480
rect 264110 -800 264222 480
rect 265292 -800 265404 480
rect 266474 -800 266586 480
rect 267656 -800 267768 480
rect 268838 -800 268950 480
rect 270020 -800 270132 480
rect 271202 -800 271314 480
rect 272384 -800 272496 480
rect 273566 -800 273678 480
rect 274748 -800 274860 480
rect 275930 -800 276042 480
rect 277112 -800 277224 480
rect 278294 -800 278406 480
rect 279476 -800 279588 480
rect 280658 -800 280770 480
rect 281840 -800 281952 480
rect 283022 -800 283134 480
rect 284204 -800 284316 480
rect 285386 -800 285498 480
rect 286568 -800 286680 480
rect 287750 -800 287862 480
rect 288932 -800 289044 480
rect 290114 -800 290226 480
rect 291296 -800 291408 480
rect 292478 -800 292590 480
rect 293660 -800 293772 480
rect 294842 -800 294954 480
rect 296024 -800 296136 480
rect 297206 -800 297318 480
rect 298388 -800 298500 480
rect 299570 -800 299682 480
rect 300752 -800 300864 480
rect 301934 -800 302046 480
rect 303116 -800 303228 480
rect 304298 -800 304410 480
rect 305480 -800 305592 480
rect 306662 -800 306774 480
rect 307844 -800 307956 480
rect 309026 -800 309138 480
rect 310208 -800 310320 480
rect 311390 -800 311502 480
rect 312572 -800 312684 480
rect 313754 -800 313866 480
rect 314936 -800 315048 480
rect 316118 -800 316230 480
rect 317300 -800 317412 480
rect 318482 -800 318594 480
rect 319664 -800 319776 480
rect 320846 -800 320958 480
rect 322028 -800 322140 480
rect 323210 -800 323322 480
rect 324392 -800 324504 480
rect 325574 -800 325686 480
rect 326756 -800 326868 480
rect 327938 -800 328050 480
rect 329120 -800 329232 480
rect 330302 -800 330414 480
rect 331484 -800 331596 480
rect 332666 -800 332778 480
rect 333848 -800 333960 480
rect 335030 -800 335142 480
rect 336212 -800 336324 480
rect 337394 -800 337506 480
rect 338576 -800 338688 480
rect 339758 -800 339870 480
rect 340940 -800 341052 480
rect 342122 -800 342234 480
rect 343304 -800 343416 480
rect 344486 -800 344598 480
rect 345668 -800 345780 480
rect 346850 -800 346962 480
rect 348032 -800 348144 480
rect 349214 -800 349326 480
rect 350396 -800 350508 480
rect 351578 -800 351690 480
rect 352760 -800 352872 480
rect 353942 -800 354054 480
rect 355124 -800 355236 480
rect 356306 -800 356418 480
rect 357488 -800 357600 480
rect 358670 -800 358782 480
rect 359852 -800 359964 480
rect 361034 -800 361146 480
rect 362216 -800 362328 480
rect 363398 -800 363510 480
rect 364580 -800 364692 480
rect 365762 -800 365874 480
rect 366944 -800 367056 480
rect 368126 -800 368238 480
rect 369308 -800 369420 480
rect 370490 -800 370602 480
rect 371672 -800 371784 480
rect 372854 -800 372966 480
rect 374036 -800 374148 480
rect 375218 -800 375330 480
rect 376400 -800 376512 480
rect 377582 -800 377694 480
rect 378764 -800 378876 480
rect 379946 -800 380058 480
rect 381128 -800 381240 480
rect 382310 -800 382422 480
rect 383492 -800 383604 480
rect 384674 -800 384786 480
rect 385856 -800 385968 480
rect 387038 -800 387150 480
rect 388220 -800 388332 480
rect 389402 -800 389514 480
rect 390584 -800 390696 480
rect 391766 -800 391878 480
rect 392948 -800 393060 480
rect 394130 -800 394242 480
rect 395312 -800 395424 480
rect 396494 -800 396606 480
rect 397676 -800 397788 480
rect 398858 -800 398970 480
rect 400040 -800 400152 480
rect 401222 -800 401334 480
rect 402404 -800 402516 480
rect 403586 -800 403698 480
rect 404768 -800 404880 480
rect 405950 -800 406062 480
rect 407132 -800 407244 480
rect 408314 -800 408426 480
rect 409496 -800 409608 480
rect 410678 -800 410790 480
rect 411860 -800 411972 480
rect 413042 -800 413154 480
rect 414224 -800 414336 480
rect 415406 -800 415518 480
rect 416588 -800 416700 480
rect 417770 -800 417882 480
rect 418952 -800 419064 480
rect 420134 -800 420246 480
rect 421316 -800 421428 480
rect 422498 -800 422610 480
rect 423680 -800 423792 480
rect 424862 -800 424974 480
rect 426044 -800 426156 480
rect 427226 -800 427338 480
rect 428408 -800 428520 480
rect 429590 -800 429702 480
rect 430772 -800 430884 480
rect 431954 -800 432066 480
rect 433136 -800 433248 480
rect 434318 -800 434430 480
rect 435500 -800 435612 480
rect 436682 -800 436794 480
rect 437864 -800 437976 480
rect 439046 -800 439158 480
rect 440228 -800 440340 480
rect 441410 -800 441522 480
rect 442592 -800 442704 480
rect 443774 -800 443886 480
rect 444956 -800 445068 480
rect 446138 -800 446250 480
rect 447320 -800 447432 480
rect 448502 -800 448614 480
rect 449684 -800 449796 480
rect 450866 -800 450978 480
rect 452048 -800 452160 480
rect 453230 -800 453342 480
rect 454412 -800 454524 480
rect 455594 -800 455706 480
rect 456776 -800 456888 480
rect 457958 -800 458070 480
rect 459140 -800 459252 480
rect 460322 -800 460434 480
rect 461504 -800 461616 480
rect 462686 -800 462798 480
rect 463868 -800 463980 480
rect 465050 -800 465162 480
rect 466232 -800 466344 480
rect 467414 -800 467526 480
rect 468596 -800 468708 480
rect 469778 -800 469890 480
rect 470960 -800 471072 480
rect 472142 -800 472254 480
rect 473324 -800 473436 480
rect 474506 -800 474618 480
rect 475688 -800 475800 480
rect 476870 -800 476982 480
rect 478052 -800 478164 480
rect 479234 -800 479346 480
rect 480416 -800 480528 480
rect 481598 -800 481710 480
rect 482780 -800 482892 480
rect 483962 -800 484074 480
rect 485144 -800 485256 480
rect 486326 -800 486438 480
rect 487508 -800 487620 480
rect 488690 -800 488802 480
rect 489872 -800 489984 480
rect 491054 -800 491166 480
rect 492236 -800 492348 480
rect 493418 -800 493530 480
rect 494600 -800 494712 480
rect 495782 -800 495894 480
rect 496964 -800 497076 480
rect 498146 -800 498258 480
rect 499328 -800 499440 480
rect 500510 -800 500622 480
rect 501692 -800 501804 480
rect 502874 -800 502986 480
rect 504056 -800 504168 480
rect 505238 -800 505350 480
rect 506420 -800 506532 480
rect 507602 -800 507714 480
rect 508784 -800 508896 480
rect 509966 -800 510078 480
rect 511148 -800 511260 480
rect 512330 -800 512442 480
rect 513512 -800 513624 480
rect 514694 -800 514806 480
rect 515876 -800 515988 480
rect 517058 -800 517170 480
rect 518240 -800 518352 480
rect 519422 -800 519534 480
rect 520604 -800 520716 480
rect 521786 -800 521898 480
rect 522968 -800 523080 480
rect 524150 -800 524262 480
rect 525332 -800 525444 480
rect 526514 -800 526626 480
rect 527696 -800 527808 480
rect 528878 -800 528990 480
rect 530060 -800 530172 480
rect 531242 -800 531354 480
rect 532424 -800 532536 480
rect 533606 -800 533718 480
rect 534788 -800 534900 480
rect 535970 -800 536082 480
rect 537152 -800 537264 480
rect 538334 -800 538446 480
rect 539516 -800 539628 480
rect 540698 -800 540810 480
rect 541880 -800 541992 480
rect 543062 -800 543174 480
rect 544244 -800 544356 480
rect 545426 -800 545538 480
rect 546608 -800 546720 480
rect 547790 -800 547902 480
rect 548972 -800 549084 480
rect 550154 -800 550266 480
rect 551336 -800 551448 480
rect 552518 -800 552630 480
rect 553700 -800 553812 480
rect 554882 -800 554994 480
rect 556064 -800 556176 480
rect 557246 -800 557358 480
rect 558428 -800 558540 480
rect 559610 -800 559722 480
rect 560792 -800 560904 480
rect 561974 -800 562086 480
rect 563156 -800 563268 480
rect 564338 -800 564450 480
rect 565520 -800 565632 480
rect 566702 -800 566814 480
rect 567884 -800 567996 480
rect 569066 -800 569178 480
rect 570248 -800 570360 480
rect 571430 -800 571542 480
rect 572612 -800 572724 480
rect 573794 -800 573906 480
rect 574976 -800 575088 480
rect 576158 -800 576270 480
rect 577340 -800 577452 480
rect 578522 -800 578634 480
rect 579704 -800 579816 480
rect 580886 -800 580998 480
rect 582068 -800 582180 480
rect 583250 -800 583362 480
<< via2 >>
rect 117052 695294 117904 695398
rect 117052 694702 117144 695294
rect 117144 694702 117816 695294
rect 117816 694702 117904 695294
rect 117052 694620 117904 694702
rect 120888 695336 122028 695502
rect 120888 694644 121002 695336
rect 121002 694644 121886 695336
rect 121886 694644 122028 695336
rect 120888 694490 122028 694644
rect 123288 695336 124428 695502
rect 123288 694644 123402 695336
rect 123402 694644 124286 695336
rect 124286 694644 124428 695336
rect 123288 694490 124428 694644
rect 127278 695396 128130 695500
rect 127278 694804 127370 695396
rect 127370 694804 128042 695396
rect 128042 694804 128130 695396
rect 127278 694722 128130 694804
rect 415460 691208 415562 691316
rect 415820 691208 415922 691316
rect 415460 690968 415562 691076
rect 415820 690968 415922 691076
rect 467360 691308 467462 691416
rect 467720 691308 467822 691416
rect 467360 691068 467462 691176
rect 467720 691068 467822 691176
rect 413812 688212 413996 688376
rect 414212 688212 414396 688376
rect 413812 687812 413996 687976
rect 414212 687812 414396 687976
rect 413812 687412 413996 687576
rect 414212 687412 414396 687576
rect 413812 687012 413996 687176
rect 414212 687012 414396 687176
rect 416212 688212 416396 688376
rect 416612 688212 416796 688376
rect 416212 687812 416396 687976
rect 416612 687812 416796 687976
rect 416212 687412 416396 687576
rect 416612 687412 416796 687576
rect 416212 687012 416396 687176
rect 416622 687012 416806 687176
rect 465812 688212 465996 688376
rect 466212 688212 466396 688376
rect 465812 687812 465996 687976
rect 466212 687812 466396 687976
rect 465812 687412 465996 687576
rect 466212 687412 466396 687576
rect 465812 687012 465996 687176
rect 466212 687012 466396 687176
rect 468212 688212 468396 688376
rect 468612 688212 468796 688376
rect 468212 687812 468396 687976
rect 468612 687812 468796 687976
rect 468212 687412 468396 687576
rect 468612 687412 468796 687576
rect 468212 687012 468396 687176
rect 468622 687012 468806 687176
rect 415460 685408 415562 685516
rect 415820 685408 415922 685516
rect 415460 685168 415562 685276
rect 415820 685168 415922 685276
rect 467360 685404 467462 685512
rect 467720 685404 467822 685512
rect 467360 685164 467462 685272
rect 467720 685164 467822 685272
rect 65052 663294 65904 663398
rect 65052 662702 65144 663294
rect 65144 662702 65816 663294
rect 65816 662702 65904 663294
rect 65052 662620 65904 662702
rect 68888 663336 70028 663502
rect 68888 662644 69002 663336
rect 69002 662644 69886 663336
rect 69886 662644 70028 663336
rect 68888 662490 70028 662644
rect 71288 663336 72428 663502
rect 71288 662644 71402 663336
rect 71402 662644 72286 663336
rect 72286 662644 72428 663336
rect 71288 662490 72428 662644
rect 75278 663396 76130 663500
rect 75278 662804 75370 663396
rect 75370 662804 76042 663396
rect 76042 662804 76130 663396
rect 75278 662722 76130 662804
rect 440260 657608 440362 657716
rect 440620 657608 440722 657716
rect 440260 657368 440362 657476
rect 440620 657368 440722 657476
rect 448860 657608 448962 657716
rect 449220 657608 449322 657716
rect 448860 657368 448962 657476
rect 449220 657368 449322 657476
rect 437812 656212 437996 656376
rect 438212 656212 438396 656376
rect 437812 655812 437996 655976
rect 438212 655812 438396 655976
rect 437812 655412 437996 655576
rect 438212 655412 438396 655576
rect 437812 655012 437996 655176
rect 438212 655012 438396 655176
rect 442412 656326 442596 656490
rect 442812 656326 442996 656490
rect 442412 655926 442596 656090
rect 442812 655926 442996 656090
rect 442412 655526 442596 655690
rect 442812 655526 442996 655690
rect 442412 655126 442596 655290
rect 442822 655126 443006 655290
rect 446212 656212 446396 656376
rect 446612 656212 446796 656376
rect 446212 655812 446396 655976
rect 446612 655812 446796 655976
rect 446212 655412 446396 655576
rect 446612 655412 446796 655576
rect 446212 655012 446396 655176
rect 446612 655012 446796 655176
rect 450812 656326 450996 656490
rect 451212 656326 451396 656490
rect 450812 655926 450996 656090
rect 451212 655926 451396 656090
rect 450812 655526 450996 655690
rect 451212 655526 451396 655690
rect 450812 655126 450996 655290
rect 451222 655126 451406 655290
rect 440260 654608 440362 654716
rect 440620 654608 440722 654716
rect 440260 654368 440362 654476
rect 440620 654368 440722 654476
rect 448860 654608 448962 654716
rect 449220 654608 449322 654716
rect 448860 654368 448962 654476
rect 449220 654368 449322 654476
rect 134560 600104 134868 600344
rect 135160 600104 135468 600344
rect 135760 600104 136068 600344
rect 136360 600104 136668 600344
rect 136960 600104 137268 600344
rect 137560 600104 137868 600344
rect 138160 600104 138468 600344
rect 134006 599540 134086 599596
rect 134126 599540 134206 599596
rect 134006 599440 134086 599496
rect 134126 599440 134206 599496
rect 140406 599540 140486 599596
rect 140526 599540 140606 599596
rect 140406 599440 140486 599496
rect 140526 599440 140606 599496
rect 134622 596998 135400 597544
rect 135822 596998 136600 597544
rect 137022 596998 137800 597544
rect 138222 596998 139000 597544
rect 85560 586104 85868 586344
rect 86160 586104 86468 586344
rect 86760 586104 87068 586344
rect 87360 586104 87668 586344
rect 87960 586104 88268 586344
rect 88560 586104 88868 586344
rect 89160 586104 89468 586344
rect 416472 586394 417092 586782
rect 438974 586180 441846 586394
rect 85006 585540 85086 585596
rect 85126 585540 85206 585596
rect 85006 585440 85086 585496
rect 85126 585440 85206 585496
rect 91406 585540 91486 585596
rect 91526 585540 91606 585596
rect 91406 585440 91486 585496
rect 91526 585440 91606 585496
rect 415878 585422 416190 585608
rect 416472 584684 417092 585072
rect 447368 584840 450242 585042
rect 85622 582998 86400 583544
rect 86822 582998 87600 583544
rect 88022 582998 88800 583544
rect 89222 582998 90000 583544
rect 101854 568504 102162 568744
rect 102454 568504 102762 568744
rect 103054 568504 103362 568744
rect 103654 568504 103962 568744
rect 104254 568504 104562 568744
rect 104854 568504 105162 568744
rect 105454 568504 105762 568744
rect 107560 568504 107868 568744
rect 108160 568504 108468 568744
rect 108760 568504 109068 568744
rect 109360 568504 109668 568744
rect 109960 568504 110268 568744
rect 110560 568504 110868 568744
rect 111160 568504 111468 568744
rect 102864 567740 102944 567796
rect 102984 567740 103064 567796
rect 102864 567640 102944 567696
rect 102984 567640 103064 567696
rect 104006 567740 104086 567796
rect 104126 567740 104206 567796
rect 104006 567640 104086 567696
rect 104126 567640 104206 567696
rect 107006 567740 107086 567796
rect 107126 567740 107206 567796
rect 107006 567640 107086 567696
rect 107126 567640 107206 567696
rect 113406 567788 113486 567844
rect 113526 567788 113606 567844
rect 113406 567688 113486 567744
rect 113526 567688 113606 567744
rect 101632 565036 102410 565582
rect 102832 565036 103610 565582
rect 104032 565036 104810 565582
rect 105232 565036 106010 565582
rect 107622 564998 108400 565544
rect 108822 564998 109600 565544
rect 110022 564998 110800 565544
rect 111222 564998 112000 565544
<< metal3 >>
rect 16194 703052 21194 704800
rect 16176 702226 21194 703052
rect 68194 702928 73194 704800
rect -800 680242 1700 685242
rect 64600 663462 66404 663994
rect 64600 662522 64982 663462
rect 65968 662522 66404 663462
rect 64600 662138 66404 662522
rect 68150 663502 73222 702928
rect 120194 702666 125194 704800
rect 120110 700232 125230 702666
rect 165594 702540 170594 704800
rect 170894 702714 173094 704800
rect 165552 702300 170594 702540
rect 170854 702300 173094 702714
rect 173394 703810 175594 704800
rect 173394 702300 175744 703810
rect 175894 702300 180894 704800
rect 217294 702300 222294 704800
rect 222594 703328 224794 704800
rect 222500 702300 224794 703328
rect 225094 702300 227294 704800
rect 227594 702300 232594 704800
rect 318994 702300 323994 704800
rect 324294 702300 326494 704800
rect 326794 702300 328994 704800
rect 329294 702300 334294 704800
rect 413394 703906 418394 704800
rect 413390 702300 418394 703906
rect 465394 702880 470394 704800
rect 510594 702892 515394 704800
rect 116600 695462 118404 695994
rect 116600 694522 116982 695462
rect 117968 694522 118404 695462
rect 116600 694138 118404 694522
rect 120128 695502 125224 700232
rect 120128 694490 120888 695502
rect 122028 694490 123288 695502
rect 124428 694490 125224 695502
rect 120128 668334 125224 694490
rect 126826 695564 128630 696096
rect 126826 694624 127208 695564
rect 128194 694624 128630 695564
rect 126826 694240 128630 694624
rect 165552 693934 170568 702300
rect 170854 692700 173082 702300
rect 170832 692140 173082 692700
rect 170832 674608 173060 692140
rect 170832 672644 173078 674608
rect 68150 662490 68888 663502
rect 70028 662490 71288 663502
rect 72428 662490 73222 663502
rect -800 643842 1660 648642
rect -800 633842 1660 638642
rect 68150 593482 73222 662490
rect 74826 663564 76630 664096
rect 74826 662624 75208 663564
rect 76194 662624 76630 663564
rect 74826 662240 76630 662624
rect 120128 657344 125218 668334
rect 170720 664214 173078 672644
rect 170584 663610 173078 664214
rect 120128 656736 125224 657344
rect 120152 652550 125224 656736
rect 170584 656290 171186 663610
rect 172478 662146 173078 663610
rect 172478 656290 172824 662146
rect 170584 655688 172824 656290
rect 67942 588042 73258 593482
rect 67914 585606 73258 588042
rect 84624 587160 90256 620620
rect 120142 617090 125286 652550
rect 173464 644306 175744 702300
rect 222500 664812 224720 702300
rect 222260 664238 224752 664812
rect 222260 656624 222764 664238
rect 224356 656624 224752 664238
rect 222260 656278 224752 656624
rect 225202 657302 227234 702300
rect 413390 691458 418372 702300
rect 465390 693606 470394 702880
rect 510580 696352 515412 702892
rect 520594 702688 525394 704800
rect 566594 702994 571594 704800
rect 520592 696352 525424 702688
rect 566592 702300 571594 702994
rect 510580 695166 525452 696352
rect 465390 693184 470416 693606
rect 465392 692464 470416 693184
rect 465390 691562 470416 692464
rect 510494 691578 525452 695166
rect 566592 694960 571574 702300
rect 546976 692176 571574 694960
rect 413376 691316 418376 691458
rect 413376 691208 415460 691316
rect 415562 691208 415820 691316
rect 415922 691208 418376 691316
rect 413376 691076 418376 691208
rect 413376 690968 415460 691076
rect 415562 690968 415820 691076
rect 415922 690968 418376 691076
rect 413376 690870 418376 690968
rect 465390 691416 470418 691562
rect 465390 691308 467360 691416
rect 467462 691308 467720 691416
rect 467822 691308 470418 691416
rect 465390 691176 470418 691308
rect 465390 691068 467360 691176
rect 467462 691068 467720 691176
rect 467822 691068 470418 691176
rect 465390 690870 470418 691068
rect 415366 690868 415684 690870
rect 466794 690864 468150 690870
rect 413730 688376 414462 688608
rect 413730 688212 413812 688376
rect 413996 688212 414212 688376
rect 414396 688212 414462 688376
rect 413730 687976 414462 688212
rect 413730 687812 413812 687976
rect 413996 687812 414212 687976
rect 414396 687812 414462 687976
rect 413730 687576 414462 687812
rect 413730 687412 413812 687576
rect 413996 687412 414212 687576
rect 414396 687412 414462 687576
rect 413730 687176 414462 687412
rect 413730 687012 413812 687176
rect 413996 687012 414212 687176
rect 414396 687012 414462 687176
rect 413730 686944 414462 687012
rect 416130 688376 416866 688598
rect 416130 688212 416212 688376
rect 416396 688212 416612 688376
rect 416796 688212 416866 688376
rect 416130 687976 416866 688212
rect 416130 687812 416212 687976
rect 416396 687812 416612 687976
rect 416796 687812 416866 687976
rect 416130 687576 416866 687812
rect 416130 687412 416212 687576
rect 416396 687412 416612 687576
rect 416796 687412 416866 687576
rect 416130 687176 416866 687412
rect 416130 687012 416212 687176
rect 416396 687012 416622 687176
rect 416806 687012 416866 687176
rect 416130 686944 416866 687012
rect 465730 688376 466466 688608
rect 465730 688212 465812 688376
rect 465996 688212 466212 688376
rect 466396 688212 466466 688376
rect 465730 687976 466466 688212
rect 465730 687812 465812 687976
rect 465996 687812 466212 687976
rect 466396 687812 466466 687976
rect 465730 687576 466466 687812
rect 465730 687412 465812 687576
rect 465996 687412 466212 687576
rect 466396 687412 466466 687576
rect 465730 687176 466466 687412
rect 465730 687012 465812 687176
rect 465996 687012 466212 687176
rect 466396 687012 466466 687176
rect 465730 686944 466466 687012
rect 468130 688376 468866 688598
rect 468130 688212 468212 688376
rect 468396 688212 468612 688376
rect 468796 688212 468866 688376
rect 468130 687976 468866 688212
rect 468130 687812 468212 687976
rect 468396 687812 468612 687976
rect 468796 687812 468866 687976
rect 468130 687576 468866 687812
rect 468130 687412 468212 687576
rect 468396 687412 468612 687576
rect 468796 687412 468866 687576
rect 468130 687176 468866 687412
rect 468130 687012 468212 687176
rect 468396 687012 468622 687176
rect 468806 687012 468866 687176
rect 468130 686944 468866 687012
rect 510494 686746 512924 691578
rect 517294 686746 519782 691578
rect 524152 687904 525452 691578
rect 524152 686746 525424 687904
rect 466650 685576 468836 685578
rect 413388 685516 418376 685576
rect 465390 685546 470376 685576
rect 413388 685408 415460 685516
rect 415562 685408 415820 685516
rect 415922 685408 418376 685516
rect 413388 685276 418376 685408
rect 413388 685168 415460 685276
rect 415562 685168 415820 685276
rect 415922 685168 418376 685276
rect 413388 684800 418376 685168
rect 465318 685512 470376 685546
rect 465318 685404 467360 685512
rect 467462 685404 467720 685512
rect 467822 685404 470376 685512
rect 465318 685272 470376 685404
rect 465318 685164 467360 685272
rect 467462 685164 467720 685272
rect 467822 685164 470376 685272
rect 465318 684800 470376 685164
rect 413390 672446 418372 684800
rect 465318 684084 470372 684800
rect 510494 684518 525424 686746
rect 465318 683036 470370 684084
rect 465318 682080 470394 683036
rect 465390 672488 470394 682080
rect 426718 672486 433774 672488
rect 426718 672446 441922 672486
rect 413390 667906 441922 672446
rect 438918 659596 441922 667906
rect 447300 667914 470394 672488
rect 447300 667900 451926 667914
rect 447318 661028 450322 667900
rect 465390 667864 470394 667914
rect 438868 657716 441950 659596
rect 447318 658442 450330 661028
rect 438868 657608 440260 657716
rect 440362 657608 440620 657716
rect 440722 657608 441950 657716
rect 438868 657476 441950 657608
rect 438868 657368 440260 657476
rect 440362 657368 440620 657476
rect 440722 657368 441950 657476
rect 225202 656220 227256 657302
rect 145408 641340 168710 641624
rect 173466 641340 175738 644306
rect 216098 641350 221908 641414
rect 225206 641350 227256 656220
rect 437730 656376 438466 656608
rect 438868 656494 441950 657368
rect 447326 657716 450330 658442
rect 447326 657608 448860 657716
rect 448962 657608 449220 657716
rect 449322 657608 450330 657716
rect 447326 657476 450330 657608
rect 447326 657368 448860 657476
rect 448962 657368 449220 657476
rect 449322 657368 450330 657476
rect 437730 656212 437812 656376
rect 437996 656212 438212 656376
rect 438396 656212 438466 656376
rect 437730 655976 438466 656212
rect 437730 655812 437812 655976
rect 437996 655812 438212 655976
rect 438396 655812 438466 655976
rect 437730 655576 438466 655812
rect 437730 655412 437812 655576
rect 437996 655412 438212 655576
rect 438396 655412 438466 655576
rect 437730 655176 438466 655412
rect 437730 655012 437812 655176
rect 437996 655012 438212 655176
rect 438396 655012 438466 655176
rect 442330 656490 443066 656712
rect 442330 656326 442412 656490
rect 442596 656326 442812 656490
rect 442996 656326 443066 656490
rect 442330 656090 443066 656326
rect 442330 655926 442412 656090
rect 442596 655926 442812 656090
rect 442996 655926 443066 656090
rect 442330 655690 443066 655926
rect 442330 655526 442412 655690
rect 442596 655526 442812 655690
rect 442996 655526 443066 655690
rect 442330 655290 443066 655526
rect 442330 655126 442412 655290
rect 442596 655126 442822 655290
rect 443006 655126 443066 655290
rect 442330 655058 443066 655126
rect 446130 656376 446866 656608
rect 447326 656540 450330 657368
rect 446130 656212 446212 656376
rect 446396 656212 446612 656376
rect 446796 656212 446866 656376
rect 446130 655976 446866 656212
rect 446130 655812 446212 655976
rect 446396 655812 446612 655976
rect 446796 655812 446866 655976
rect 446130 655576 446866 655812
rect 446130 655412 446212 655576
rect 446396 655412 446612 655576
rect 446796 655412 446866 655576
rect 446130 655176 446866 655412
rect 437730 654944 438466 655012
rect 438924 655022 441930 655024
rect 438924 654716 441974 655022
rect 446130 655012 446212 655176
rect 446396 655012 446612 655176
rect 446796 655012 446866 655176
rect 450730 656490 451466 656712
rect 450730 656326 450812 656490
rect 450996 656326 451212 656490
rect 451396 656326 451466 656490
rect 450730 656090 451466 656326
rect 450730 655926 450812 656090
rect 450996 655926 451212 656090
rect 451396 655926 451466 656090
rect 450730 655690 451466 655926
rect 450730 655526 450812 655690
rect 450996 655526 451212 655690
rect 451396 655526 451466 655690
rect 450730 655290 451466 655526
rect 450730 655126 450812 655290
rect 450996 655126 451222 655290
rect 451406 655126 451466 655290
rect 450730 655058 451466 655126
rect 446130 654944 446866 655012
rect 438924 654608 440260 654716
rect 440362 654608 440620 654716
rect 440722 654714 441974 654716
rect 447300 654716 450342 654936
rect 440722 654608 441968 654714
rect 438924 654476 441968 654608
rect 438924 654368 440260 654476
rect 440362 654368 440620 654476
rect 440722 654368 441968 654476
rect 438924 651142 441968 654368
rect 447300 654608 448860 654716
rect 448962 654608 449220 654716
rect 449322 654608 450342 654716
rect 447300 654476 450342 654608
rect 447300 654368 448860 654476
rect 448962 654368 449220 654476
rect 449322 654368 450342 654476
rect 447300 653986 450342 654368
rect 438918 650114 441968 651142
rect 447316 651142 450320 653986
rect 227664 641350 238982 641414
rect 145408 641306 170068 641340
rect 173362 641316 179734 641340
rect 216098 641316 238982 641350
rect 351700 641316 362636 641330
rect 145408 641300 172954 641306
rect 173362 641300 362636 641316
rect 145408 639526 362636 641300
rect 145408 633438 354208 639526
rect 360382 633438 362636 639526
rect 145408 631824 362636 633438
rect 145408 631774 294570 631824
rect 145408 631608 168710 631774
rect 177012 631742 294570 631774
rect 216098 631660 238982 631742
rect 120152 610410 125224 617090
rect 120120 608504 125224 610410
rect 120120 600802 125138 608504
rect 133624 601160 139256 603044
rect 120132 599628 125126 600802
rect 133620 600344 139258 601160
rect 133620 600104 134560 600344
rect 134868 600104 135160 600344
rect 135468 600104 135760 600344
rect 136068 600104 136360 600344
rect 136668 600104 136960 600344
rect 137268 600104 137560 600344
rect 137868 600104 138160 600344
rect 138468 600104 139258 600344
rect 133620 600020 139258 600104
rect 145042 599640 145378 599646
rect 120132 599606 132244 599628
rect 142080 599606 145378 599640
rect 120132 599596 134274 599606
rect 120132 599540 134006 599596
rect 134086 599540 134126 599596
rect 134206 599540 134274 599596
rect 120132 599496 134274 599540
rect 120132 599440 134006 599496
rect 134086 599440 134126 599496
rect 134206 599440 134274 599496
rect 120132 599412 134274 599440
rect 140370 599596 145378 599606
rect 140370 599540 140406 599596
rect 140486 599540 140526 599596
rect 140606 599540 145378 599596
rect 140370 599496 145378 599540
rect 140370 599440 140406 599496
rect 140486 599440 140526 599496
rect 140606 599440 145378 599496
rect 140370 599412 145378 599440
rect 120132 599370 132244 599412
rect 133984 599410 134258 599412
rect 140384 599410 140628 599412
rect 142080 599394 145378 599412
rect 120132 599278 125126 599370
rect 134234 597544 139146 597958
rect 134234 596998 134622 597544
rect 135400 596998 135822 597544
rect 136600 596998 137022 597544
rect 137800 596998 138222 597544
rect 139000 596998 139146 597544
rect 134234 596602 139146 596998
rect 145042 587836 145378 599394
rect 208174 587836 211476 587926
rect 145042 587620 421640 587836
rect 145042 587562 145378 587620
rect 208174 587372 211476 587620
rect 84620 586344 90258 587160
rect 421178 587112 421598 587620
rect 84620 586104 85560 586344
rect 85868 586104 86160 586344
rect 86468 586104 86760 586344
rect 87068 586104 87360 586344
rect 87668 586104 87960 586344
rect 88268 586104 88560 586344
rect 88868 586104 89160 586344
rect 89468 586104 90258 586344
rect 416354 586782 417192 586912
rect 416354 586394 416472 586782
rect 417092 586394 417192 586782
rect 416354 586296 417192 586394
rect 438918 586394 441922 650114
rect 447316 649884 450322 651142
rect 447318 586662 450322 649884
rect 547102 632150 550106 692176
rect 566592 692132 571574 692176
rect 582300 677984 584800 682984
rect 565206 644596 576142 646006
rect 565206 644584 583128 644596
rect 565206 644560 584800 644584
rect 565206 641590 567706 644560
rect 564368 639756 567706 641590
rect 573760 639812 584800 644560
rect 573760 639756 576142 639812
rect 582340 639784 584800 639812
rect 564368 634590 576142 639756
rect 564368 634584 583082 634590
rect 564368 634562 584800 634584
rect 547102 629150 550128 632150
rect 564368 632060 567668 634562
rect 447316 586398 450322 586662
rect 438918 586356 438974 586394
rect 84620 586020 90258 586104
rect 438908 586180 438974 586356
rect 441846 586356 441922 586394
rect 441846 586180 441924 586356
rect 438908 586102 441924 586180
rect 447312 586048 450322 586398
rect 127102 585626 129270 585630
rect 115776 585620 129270 585626
rect 104672 585606 129270 585620
rect 415786 585614 416282 585710
rect 415786 585608 417586 585614
rect 415786 585606 415878 585608
rect 67914 585596 85274 585606
rect 67914 585540 85006 585596
rect 85086 585540 85126 585596
rect 85206 585540 85274 585596
rect 67914 585496 85274 585540
rect 67914 585440 85006 585496
rect 85086 585440 85126 585496
rect 85206 585440 85274 585496
rect 67914 585412 85274 585440
rect 91370 585604 218504 585606
rect 230148 585604 402784 585606
rect 91370 585600 402784 585604
rect 412402 585600 415878 585606
rect 91370 585596 415878 585600
rect 91370 585540 91406 585596
rect 91486 585540 91526 585596
rect 91606 585540 415878 585596
rect 91370 585496 415878 585540
rect 91370 585440 91406 585496
rect 91486 585440 91526 585496
rect 91606 585440 415878 585496
rect 91370 585422 415878 585440
rect 416190 585422 417586 585608
rect 91370 585412 417586 585422
rect 447316 585414 450318 586048
rect 67914 585282 73258 585412
rect 84984 585410 85258 585412
rect 91384 585410 91628 585412
rect 104672 585386 129270 585412
rect 218288 585410 230804 585412
rect 402662 585406 412608 585412
rect 104672 585380 116174 585386
rect 118856 585382 122066 585386
rect 127102 585374 129270 585386
rect 415786 585344 416282 585412
rect 67914 567806 73226 585282
rect 447312 585258 450318 585414
rect 416354 585072 417186 585172
rect 416354 584684 416472 585072
rect 417092 584684 417186 585072
rect 447312 585042 450316 585258
rect 447312 584840 447368 585042
rect 450242 584840 450316 585042
rect 447312 584780 450316 584840
rect 416354 584586 417186 584684
rect 85234 583544 90146 583958
rect 85234 582998 85622 583544
rect 86400 582998 86822 583544
rect 87600 582998 88022 583544
rect 88800 582998 89222 583544
rect 90000 582998 90146 583544
rect 85234 582602 90146 582998
rect 101388 568744 106034 569082
rect 101388 568504 101854 568744
rect 102162 568504 102454 568744
rect 102762 568504 103054 568744
rect 103362 568504 103654 568744
rect 103962 568504 104254 568744
rect 104562 568504 104854 568744
rect 105162 568504 105454 568744
rect 105762 568504 106034 568744
rect 101388 568420 106034 568504
rect 107094 568744 111740 569082
rect 107094 568504 107560 568744
rect 107868 568504 108160 568744
rect 108468 568504 108760 568744
rect 109068 568504 109360 568744
rect 109668 568504 109960 568744
rect 110268 568504 110560 568744
rect 110868 568504 111160 568744
rect 111468 568504 111740 568744
rect 107094 568420 111740 568504
rect 116646 567854 124748 567860
rect 547124 567854 550128 629150
rect 565206 629758 567668 632060
rect 573722 629784 584800 634562
rect 573722 629758 576142 629784
rect 565206 627532 576142 629758
rect 583520 589472 584800 589584
rect 583520 588290 584800 588402
rect 583520 587108 584800 587220
rect 583520 585926 584800 586038
rect 583520 584744 584800 584856
rect 583520 583562 584800 583674
rect 113382 567844 550128 567854
rect 102338 567806 102860 567808
rect 67914 567796 103076 567806
rect 67914 567740 102864 567796
rect 102944 567740 102984 567796
rect 103064 567740 103076 567796
rect 67914 567696 103076 567740
rect 67914 567640 102864 567696
rect 102944 567640 102984 567696
rect 103064 567640 103076 567696
rect 67914 567610 103076 567640
rect 103986 567796 107220 567806
rect 103986 567740 104006 567796
rect 104086 567740 104126 567796
rect 104206 567740 107006 567796
rect 107086 567740 107126 567796
rect 107206 567740 107220 567796
rect 103986 567696 107220 567740
rect 103986 567640 104006 567696
rect 104086 567640 104126 567696
rect 104206 567640 107006 567696
rect 107086 567640 107126 567696
rect 107206 567640 107220 567696
rect 113382 567788 113406 567844
rect 113486 567788 113526 567844
rect 113606 567788 550128 567844
rect 113382 567744 550128 567788
rect 113382 567688 113406 567744
rect 113486 567688 113526 567744
rect 113606 567688 550128 567744
rect 113382 567658 550128 567688
rect 113472 567654 113606 567658
rect 116646 567640 124748 567658
rect 547124 567642 550128 567658
rect 103986 567610 107220 567640
rect 67914 567600 73226 567610
rect 102338 567606 102860 567610
rect 101244 565582 106156 565996
rect 101244 565036 101632 565582
rect 102410 565036 102832 565582
rect 103610 565036 104032 565582
rect 104810 565036 105232 565582
rect 106010 565036 106156 565582
rect 101244 564640 106156 565036
rect 107234 565544 112146 565958
rect 107234 564998 107622 565544
rect 108400 564998 108822 565544
rect 109600 564998 110022 565544
rect 110800 564998 111222 565544
rect 112000 564998 112146 565544
rect 107234 564602 112146 564998
rect -800 559442 1660 564242
rect -800 549442 1660 554242
rect 582340 550562 584800 555362
rect 582340 540562 584800 545362
rect -800 511530 480 511642
rect -800 510348 480 510460
rect -800 509166 480 509278
rect -800 507984 480 508096
rect -800 506802 480 506914
rect -800 505620 480 505732
rect 583520 500050 584800 500162
rect 583520 498868 584800 498980
rect 583520 497686 584800 497798
rect 583520 496504 584800 496616
rect 583520 495322 584800 495434
rect 583520 494140 584800 494252
rect -800 468308 480 468420
rect -800 467126 480 467238
rect -800 465944 480 466056
rect -800 464762 480 464874
rect -800 463580 480 463692
rect -800 462398 480 462510
rect 583520 455628 584800 455740
rect 583520 454446 584800 454558
rect 583520 453264 584800 453376
rect 583520 452082 584800 452194
rect 583520 450900 584800 451012
rect 583520 449718 584800 449830
rect -800 425086 480 425198
rect -800 423904 480 424016
rect -800 422722 480 422834
rect -800 421540 480 421652
rect -800 420358 480 420470
rect -800 419176 480 419288
rect 583520 411206 584800 411318
rect 583520 410024 584800 410136
rect 583520 408842 584800 408954
rect 583520 407660 584800 407772
rect 583520 406478 584800 406590
rect 583520 405296 584800 405408
rect -800 381864 480 381976
rect -800 380682 480 380794
rect -800 379500 480 379612
rect -800 378318 480 378430
rect -800 377136 480 377248
rect -800 375954 480 376066
rect 583520 364784 584800 364896
rect 583520 363602 584800 363714
rect 583520 362420 584800 362532
rect 583520 361238 584800 361350
rect 583520 360056 584800 360168
rect 583520 358874 584800 358986
rect -800 338642 480 338754
rect -800 337460 480 337572
rect -800 336278 480 336390
rect -800 335096 480 335208
rect -800 333914 480 334026
rect -800 332732 480 332844
rect 583520 319562 584800 319674
rect 583520 318380 584800 318492
rect 583520 317198 584800 317310
rect 583520 316016 584800 316128
rect 583520 314834 584800 314946
rect 583520 313652 584800 313764
rect -800 295420 480 295532
rect -800 294238 480 294350
rect -800 293056 480 293168
rect -800 291874 480 291986
rect -800 290692 480 290804
rect -800 289510 480 289622
rect 583520 275140 584800 275252
rect 583520 273958 584800 274070
rect 583520 272776 584800 272888
rect 583520 271594 584800 271706
rect 583520 270412 584800 270524
rect 583520 269230 584800 269342
rect -800 252398 480 252510
rect -800 251216 480 251328
rect -800 250034 480 250146
rect -800 248852 480 248964
rect -800 247670 480 247782
rect -800 246488 480 246600
rect 582340 235230 584800 240030
rect 582340 225230 584800 230030
rect -800 214888 1660 219688
rect -800 204888 1660 209688
rect 582188 196230 582876 196238
rect 582188 191430 584800 196230
rect 582188 191424 582876 191430
rect 582340 186224 584800 186230
rect 582188 181430 584800 186224
rect 582188 181410 582678 181430
rect -800 172888 1660 177688
rect -800 162888 1660 167688
rect 582340 151538 584800 151630
rect 581994 146830 584800 151538
rect 581994 146778 583364 146830
rect 581994 141630 583088 141672
rect 581994 136912 584800 141630
rect 582340 136830 584800 136912
rect -800 124776 480 124888
rect -800 123594 480 123706
rect -800 122412 480 122524
rect -800 121230 480 121342
rect -800 120048 480 120160
rect -800 118866 480 118978
rect 583520 95118 584800 95230
rect 583520 93936 584800 94048
rect 583520 92754 584800 92866
rect 583520 91572 584800 91684
rect -800 81554 480 81666
rect -800 80372 480 80484
rect -800 79190 480 79302
rect -800 78008 480 78120
rect -800 76826 480 76938
rect -800 75644 480 75756
rect 583520 50460 584800 50572
rect 583520 49278 584800 49390
rect 583520 48096 584800 48208
rect 583520 46914 584800 47026
rect -800 38332 480 38444
rect -800 37150 480 37262
rect -800 35968 480 36080
rect -800 34786 480 34898
rect -800 33604 480 33716
rect -800 32422 480 32534
rect 583520 24002 584800 24114
rect 583520 22820 584800 22932
rect 583520 21638 584800 21750
rect 583520 20456 584800 20568
rect 583520 19274 584800 19386
rect 583520 18092 584800 18204
rect -800 16910 480 17022
rect 583520 16910 584800 17022
rect -800 15728 480 15840
rect 583520 15728 584800 15840
rect -800 14546 480 14658
rect 583520 14546 584800 14658
rect -800 13364 480 13476
rect 583520 13364 584800 13476
rect -800 12182 480 12294
rect 583520 12182 584800 12294
rect -800 11000 480 11112
rect 583520 11000 584800 11112
rect -800 9818 480 9930
rect 583520 9818 584800 9930
rect -800 8636 480 8748
rect 583520 8636 584800 8748
rect -800 7454 480 7566
rect 583520 7454 584800 7566
rect -800 6272 480 6384
rect 583520 6272 584800 6384
rect -800 5090 480 5202
rect 583520 5090 584800 5202
rect -800 3908 480 4020
rect 583520 3908 584800 4020
rect -800 2726 480 2838
rect 583520 2726 584800 2838
rect -800 1544 480 1656
rect 583520 1544 584800 1656
<< via3 >>
rect 64982 663398 65968 663462
rect 64982 662620 65052 663398
rect 65052 662620 65904 663398
rect 65904 662620 65968 663398
rect 64982 662522 65968 662620
rect 116982 695398 117968 695462
rect 116982 694620 117052 695398
rect 117052 694620 117904 695398
rect 117904 694620 117968 695398
rect 116982 694522 117968 694620
rect 127208 695500 128194 695564
rect 127208 694722 127278 695500
rect 127278 694722 128130 695500
rect 128130 694722 128194 695500
rect 127208 694624 128194 694722
rect 75208 663500 76194 663564
rect 75208 662722 75278 663500
rect 75278 662722 76130 663500
rect 76130 662722 76194 663500
rect 75208 662624 76194 662722
rect 171186 656290 172478 663610
rect 222764 656624 224356 664238
rect 413812 688212 413996 688376
rect 414212 688212 414396 688376
rect 413812 687812 413996 687976
rect 414212 687812 414396 687976
rect 413812 687412 413996 687576
rect 414212 687412 414396 687576
rect 413812 687012 413996 687176
rect 414212 687012 414396 687176
rect 416212 688212 416396 688376
rect 416612 688212 416796 688376
rect 416212 687812 416396 687976
rect 416612 687812 416796 687976
rect 416212 687412 416396 687576
rect 416612 687412 416796 687576
rect 416212 687012 416396 687176
rect 416622 687012 416806 687176
rect 465812 688212 465996 688376
rect 466212 688212 466396 688376
rect 465812 687812 465996 687976
rect 466212 687812 466396 687976
rect 465812 687412 465996 687576
rect 466212 687412 466396 687576
rect 465812 687012 465996 687176
rect 466212 687012 466396 687176
rect 468212 688212 468396 688376
rect 468612 688212 468796 688376
rect 468212 687812 468396 687976
rect 468612 687812 468796 687976
rect 468212 687412 468396 687576
rect 468612 687412 468796 687576
rect 468212 687012 468396 687176
rect 468622 687012 468806 687176
rect 512924 686746 517294 691578
rect 519782 686746 524152 691578
rect 437812 656212 437996 656376
rect 438212 656212 438396 656376
rect 437812 655812 437996 655976
rect 438212 655812 438396 655976
rect 437812 655412 437996 655576
rect 438212 655412 438396 655576
rect 437812 655012 437996 655176
rect 438212 655012 438396 655176
rect 442412 656326 442596 656490
rect 442812 656326 442996 656490
rect 442412 655926 442596 656090
rect 442812 655926 442996 656090
rect 442412 655526 442596 655690
rect 442812 655526 442996 655690
rect 442412 655126 442596 655290
rect 442822 655126 443006 655290
rect 446212 656212 446396 656376
rect 446612 656212 446796 656376
rect 446212 655812 446396 655976
rect 446612 655812 446796 655976
rect 446212 655412 446396 655576
rect 446612 655412 446796 655576
rect 446212 655012 446396 655176
rect 446612 655012 446796 655176
rect 450812 656326 450996 656490
rect 451212 656326 451396 656490
rect 450812 655926 450996 656090
rect 451212 655926 451396 656090
rect 450812 655526 450996 655690
rect 451212 655526 451396 655690
rect 450812 655126 450996 655290
rect 451222 655126 451406 655290
rect 354208 633438 360382 639526
rect 134560 600104 134868 600344
rect 135160 600104 135468 600344
rect 135760 600104 136068 600344
rect 136360 600104 136668 600344
rect 136960 600104 137268 600344
rect 137560 600104 137868 600344
rect 138160 600104 138468 600344
rect 134622 596998 135400 597544
rect 135822 596998 136600 597544
rect 137022 596998 137800 597544
rect 138222 596998 139000 597544
rect 85560 586104 85868 586344
rect 86160 586104 86468 586344
rect 86760 586104 87068 586344
rect 87360 586104 87668 586344
rect 87960 586104 88268 586344
rect 88560 586104 88868 586344
rect 89160 586104 89468 586344
rect 416472 586394 417092 586782
rect 567706 639756 573760 644560
rect 416472 584684 417092 585072
rect 85622 582998 86400 583544
rect 86822 582998 87600 583544
rect 88022 582998 88800 583544
rect 89222 582998 90000 583544
rect 101854 568504 102162 568744
rect 102454 568504 102762 568744
rect 103054 568504 103362 568744
rect 103654 568504 103962 568744
rect 104254 568504 104562 568744
rect 104854 568504 105162 568744
rect 105454 568504 105762 568744
rect 107560 568504 107868 568744
rect 108160 568504 108468 568744
rect 108760 568504 109068 568744
rect 109360 568504 109668 568744
rect 109960 568504 110268 568744
rect 110560 568504 110868 568744
rect 111160 568504 111468 568744
rect 567668 629758 573722 634562
rect 101632 565036 102410 565582
rect 102832 565036 103610 565582
rect 104032 565036 104810 565582
rect 105232 565036 106010 565582
rect 107622 564998 108400 565544
rect 108822 564998 109600 565544
rect 110022 564998 110800 565544
rect 111222 564998 112000 565544
<< metal4 >>
rect 165594 702540 170594 704800
rect 141374 696222 153568 702508
rect 128194 696172 153568 696222
rect 116600 695542 118404 695994
rect 116600 694458 116918 695542
rect 118020 694458 118404 695542
rect 116600 694138 118404 694458
rect 126746 695564 153568 696172
rect 126746 694624 127208 695564
rect 128194 694624 153568 695564
rect 126746 694244 153568 694624
rect 126826 694240 128630 694244
rect 74746 664108 78146 664172
rect 84288 664108 96474 681736
rect 141374 681172 153568 694244
rect 165552 702300 170594 702540
rect 175894 702434 180894 704800
rect 175862 702300 180894 702434
rect 217294 702970 222294 704800
rect 217294 702300 222336 702970
rect 227594 702926 232594 704800
rect 165552 696162 170568 702300
rect 165552 693934 170584 696162
rect 165554 682686 170584 693934
rect 175862 682686 180868 702300
rect 217306 684124 222336 702300
rect 165508 682660 187874 682686
rect 217280 682660 222336 684124
rect 227582 694624 232594 702926
rect 318994 702300 323994 704800
rect 329294 702300 334294 704800
rect 227582 682660 232548 694624
rect 402706 694056 476700 696958
rect 402738 688608 404890 694056
rect 412670 688608 414760 688612
rect 463316 688610 464766 694056
rect 511622 691578 524816 694356
rect 402692 688376 414760 688608
rect 463308 688608 465444 688610
rect 416124 688598 416882 688604
rect 402692 688212 413812 688376
rect 413996 688212 414212 688376
rect 414396 688212 414760 688376
rect 402692 687976 414760 688212
rect 402692 687812 413812 687976
rect 413996 687812 414212 687976
rect 414396 687812 414760 687976
rect 402692 687576 414760 687812
rect 402692 687412 413812 687576
rect 413996 687412 414212 687576
rect 414396 687412 414760 687576
rect 402692 687176 414760 687412
rect 402692 687012 413812 687176
rect 413996 687012 414212 687176
rect 414396 687012 414760 687176
rect 402692 686948 414760 687012
rect 416120 688376 416882 688598
rect 416120 688212 416212 688376
rect 416396 688212 416612 688376
rect 416796 688212 416882 688376
rect 416120 688050 416882 688212
rect 416120 688042 416560 688050
rect 416120 687738 416166 688042
rect 416450 687746 416560 688042
rect 416844 687746 416882 688050
rect 416450 687738 416882 687746
rect 416120 687576 416882 687738
rect 416120 687412 416212 687576
rect 416396 687412 416612 687576
rect 416796 687412 416882 687576
rect 416120 687258 416882 687412
rect 416120 686962 416156 687258
rect 416484 687254 416882 687258
rect 416484 686962 416568 687254
rect 416120 686950 416568 686962
rect 416852 686950 416882 687254
rect 416120 686948 416882 686950
rect 165508 682658 191410 682660
rect 208250 682658 232548 682660
rect 64600 663542 66404 663994
rect 64600 662458 64918 663542
rect 66020 662458 66404 663542
rect 64600 662138 66404 662458
rect 74746 663564 96474 664108
rect 74746 662624 75208 663564
rect 76194 662624 96474 663564
rect 74746 662262 96474 662624
rect 74746 662244 78146 662262
rect 74826 662240 76630 662244
rect 84288 641240 96474 662262
rect 141380 641240 153566 681172
rect 165508 677212 191570 682658
rect 185918 677168 191570 677212
rect 186722 676918 191570 677168
rect 204138 677168 232548 682658
rect 402730 681322 404890 686948
rect 412670 686942 414760 686948
rect 416124 686946 416882 686948
rect 463308 688376 466460 688608
rect 468124 688598 468882 688604
rect 463308 688212 465812 688376
rect 465996 688212 466212 688376
rect 466396 688212 466460 688376
rect 463308 687976 466460 688212
rect 463308 687812 465812 687976
rect 465996 687812 466212 687976
rect 466396 687812 466460 687976
rect 463308 687576 466460 687812
rect 463308 687412 465812 687576
rect 465996 687412 466212 687576
rect 466396 687412 466460 687576
rect 463308 687176 466460 687412
rect 463308 687012 465812 687176
rect 465996 687012 466212 687176
rect 466396 687012 466460 687176
rect 463308 686948 466460 687012
rect 468120 688376 468882 688598
rect 468120 688212 468212 688376
rect 468396 688212 468612 688376
rect 468796 688212 468882 688376
rect 468120 688050 468882 688212
rect 468120 688042 468560 688050
rect 468120 687738 468166 688042
rect 468450 687746 468560 688042
rect 468844 687746 468882 688050
rect 468450 687738 468882 687746
rect 468120 687576 468882 687738
rect 468120 687412 468212 687576
rect 468396 687412 468612 687576
rect 468796 687412 468882 687576
rect 468120 687258 468882 687412
rect 468120 686962 468156 687258
rect 468484 687254 468882 687258
rect 468484 686962 468568 687254
rect 468120 686950 468568 686962
rect 468852 686950 468882 687254
rect 468120 686948 468882 686950
rect 463308 686946 465444 686948
rect 468124 686946 468882 686948
rect 511622 686746 512924 691578
rect 517294 686746 519782 691578
rect 524152 686746 524816 691578
rect 511622 684546 524816 686746
rect 204138 676918 209704 677168
rect 222268 664238 224752 664696
rect 170584 663610 172824 664214
rect 170584 656290 171186 663610
rect 172478 661626 172824 663610
rect 222268 661626 222764 664238
rect 172478 661560 185306 661626
rect 213460 661560 222764 661626
rect 172478 658966 222764 661560
rect 172478 656290 172824 658966
rect 181400 658866 215482 658966
rect 170584 655688 172824 656290
rect 222268 656624 222764 658966
rect 224356 656624 224752 664238
rect 222268 656278 224752 656624
rect 402730 641404 404778 681322
rect 442324 656712 443082 656718
rect 450724 656712 451482 656718
rect 437706 656562 438460 656608
rect 434474 656552 438460 656562
rect 431788 656376 438460 656552
rect 431788 656212 437812 656376
rect 437996 656212 438212 656376
rect 438396 656212 438460 656376
rect 431788 655976 438460 656212
rect 431788 655812 437812 655976
rect 437996 655812 438212 655976
rect 438396 655812 438460 655976
rect 431788 655576 438460 655812
rect 431788 655412 437812 655576
rect 437996 655412 438212 655576
rect 438396 655412 438460 655576
rect 431788 655176 438460 655412
rect 431788 655012 437812 655176
rect 437996 655012 438212 655176
rect 438396 655012 438460 655176
rect 442320 656490 443082 656712
rect 446106 656562 446860 656608
rect 445486 656560 446860 656562
rect 442320 656326 442412 656490
rect 442596 656326 442812 656490
rect 442996 656326 443082 656490
rect 442320 656164 443082 656326
rect 442320 656156 442760 656164
rect 442320 655852 442366 656156
rect 442650 655860 442760 656156
rect 443044 655860 443082 656164
rect 442650 655852 443082 655860
rect 442320 655690 443082 655852
rect 442320 655526 442412 655690
rect 442596 655526 442812 655690
rect 442996 655526 443082 655690
rect 442320 655372 443082 655526
rect 442320 655076 442356 655372
rect 442684 655368 443082 655372
rect 442684 655076 442768 655368
rect 442320 655064 442768 655076
rect 443052 655064 443082 655368
rect 442320 655062 443082 655064
rect 442324 655060 443082 655062
rect 443936 656376 446860 656560
rect 443936 656212 446212 656376
rect 446396 656212 446612 656376
rect 446796 656212 446860 656376
rect 443936 655976 446860 656212
rect 443936 655812 446212 655976
rect 446396 655812 446612 655976
rect 446796 655812 446860 655976
rect 443936 655576 446860 655812
rect 443936 655412 446212 655576
rect 446396 655412 446612 655576
rect 446796 655412 446860 655576
rect 443936 655176 446860 655412
rect 431788 654976 438460 655012
rect 431788 641404 433780 654976
rect 437706 654948 438460 654976
rect 443936 655012 446212 655176
rect 446396 655012 446612 655176
rect 446796 655012 446860 655176
rect 450720 656490 451482 656712
rect 450720 656326 450812 656490
rect 450996 656326 451212 656490
rect 451396 656326 451482 656490
rect 450720 656164 451482 656326
rect 450720 656156 451160 656164
rect 450720 655852 450766 656156
rect 451050 655860 451160 656156
rect 451444 655860 451482 656164
rect 451050 655852 451482 655860
rect 450720 655690 451482 655852
rect 450720 655526 450812 655690
rect 450996 655526 451212 655690
rect 451396 655526 451482 655690
rect 450720 655372 451482 655526
rect 450720 655076 450756 655372
rect 451084 655368 451482 655372
rect 451084 655076 451168 655368
rect 450720 655064 451168 655076
rect 451452 655064 451482 655368
rect 450720 655062 451482 655064
rect 450724 655060 451482 655062
rect 443936 654976 446860 655012
rect 443936 641404 445822 654976
rect 446106 654948 446860 654976
rect 565206 644560 576142 646006
rect 565206 641590 567706 644560
rect 476622 641404 567706 641590
rect 351700 641284 362636 641330
rect 400454 641284 567706 641404
rect 351700 641240 567706 641284
rect 84288 639756 567706 641240
rect 573760 639756 576142 644560
rect 84288 639526 576142 639756
rect 84288 633438 354208 639526
rect 360382 634562 576142 639526
rect 360382 633438 567668 634562
rect 84288 632060 567668 633438
rect 84288 631874 495080 632060
rect 84288 631824 374398 631874
rect 402730 631868 404778 631874
rect 84288 630674 294570 631824
rect 84288 630456 96474 630674
rect 84472 586344 90336 630456
rect 84472 586130 85560 586344
rect 85148 586104 85560 586130
rect 85868 586104 86160 586344
rect 86468 586104 86760 586344
rect 87068 586104 87360 586344
rect 87668 586104 87960 586344
rect 88268 586104 88560 586344
rect 88868 586104 89160 586344
rect 89468 586130 90336 586344
rect 101248 587156 111738 630674
rect 133558 603044 139362 630674
rect 186722 630654 191570 630674
rect 204138 630654 209704 630674
rect 133472 602336 139362 603044
rect 133472 600344 139336 602336
rect 133472 600130 134560 600344
rect 134148 600104 134560 600130
rect 134868 600104 135160 600344
rect 135468 600104 135760 600344
rect 136068 600104 136360 600344
rect 136668 600104 136960 600344
rect 137268 600104 137560 600344
rect 137868 600104 138160 600344
rect 138468 600130 139336 600344
rect 138468 600104 139080 600130
rect 134148 600024 139080 600104
rect 134148 600014 134494 600024
rect 134234 597544 139146 597958
rect 134234 596998 134622 597544
rect 135400 596998 135822 597544
rect 136600 596998 137022 597544
rect 137800 596998 138222 597544
rect 139000 596998 139146 597544
rect 134234 596602 139146 596998
rect 417434 591470 424178 631874
rect 565206 629758 567668 632060
rect 573722 629758 576142 634562
rect 565206 627532 576142 629758
rect 417438 590348 424178 591470
rect 417438 589372 424184 590348
rect 417438 588084 424158 589372
rect 89468 586104 90080 586130
rect 85148 586024 90080 586104
rect 85148 586014 85494 586024
rect 85234 583544 90146 583958
rect 85234 582998 85622 583544
rect 86400 582998 86822 583544
rect 87600 582998 88022 583544
rect 88800 582998 89222 583544
rect 90000 582998 90146 583544
rect 85234 582602 90146 582998
rect 101248 582374 111700 587156
rect 416354 586782 417192 586912
rect 416354 586394 416472 586782
rect 417092 586394 417192 586782
rect 416354 586296 417192 586394
rect 416354 585072 417186 585172
rect 416354 584684 416472 585072
rect 417092 584684 417186 585072
rect 416354 584586 417186 584684
rect 101248 577176 111738 582374
rect 101404 570812 111738 577176
rect 101374 569594 111738 570812
rect 101386 569170 111738 569594
rect 101388 568854 111738 569170
rect 101388 568744 111740 568854
rect 101388 568504 101854 568744
rect 102162 568504 102454 568744
rect 102762 568504 103054 568744
rect 103362 568504 103654 568744
rect 103962 568504 104254 568744
rect 104562 568504 104854 568744
rect 105162 568504 105454 568744
rect 105762 568504 107560 568744
rect 107868 568504 108160 568744
rect 108468 568504 108760 568744
rect 109068 568504 109360 568744
rect 109668 568504 109960 568744
rect 110268 568504 110560 568744
rect 110868 568504 111160 568744
rect 111468 568504 111740 568744
rect 101388 568424 111740 568504
rect 101388 568414 101788 568424
rect 105804 568420 107494 568424
rect 107094 568414 107494 568420
rect 101244 565582 106156 565996
rect 101244 565036 101632 565582
rect 102410 565036 102832 565582
rect 103610 565036 104032 565582
rect 104810 565036 105232 565582
rect 106010 565036 106156 565582
rect 101244 564640 106156 565036
rect 107234 565544 112146 565958
rect 107234 564998 107622 565544
rect 108400 564998 108822 565544
rect 109600 564998 110022 565544
rect 110800 564998 111222 565544
rect 112000 564998 112146 565544
rect 107234 564602 112146 564998
<< via4 >>
rect 116918 695462 118020 695542
rect 116918 694522 116982 695462
rect 116982 694522 117968 695462
rect 117968 694522 118020 695462
rect 116918 694458 118020 694522
rect 416166 687976 416450 688042
rect 416166 687812 416212 687976
rect 416212 687812 416396 687976
rect 416396 687812 416450 687976
rect 416166 687738 416450 687812
rect 416560 687976 416844 688050
rect 416560 687812 416612 687976
rect 416612 687812 416796 687976
rect 416796 687812 416844 687976
rect 416560 687746 416844 687812
rect 416156 687176 416484 687258
rect 416156 687012 416212 687176
rect 416212 687012 416396 687176
rect 416396 687012 416484 687176
rect 416156 686962 416484 687012
rect 416568 687176 416852 687254
rect 416568 687012 416622 687176
rect 416622 687012 416806 687176
rect 416806 687012 416852 687176
rect 416568 686950 416852 687012
rect 64918 663462 66020 663542
rect 64918 662522 64982 663462
rect 64982 662522 65968 663462
rect 65968 662522 66020 663462
rect 64918 662458 66020 662522
rect 468166 687976 468450 688042
rect 468166 687812 468212 687976
rect 468212 687812 468396 687976
rect 468396 687812 468450 687976
rect 468166 687738 468450 687812
rect 468560 687976 468844 688050
rect 468560 687812 468612 687976
rect 468612 687812 468796 687976
rect 468796 687812 468844 687976
rect 468560 687746 468844 687812
rect 468156 687176 468484 687258
rect 468156 687012 468212 687176
rect 468212 687012 468396 687176
rect 468396 687012 468484 687176
rect 468156 686962 468484 687012
rect 468568 687176 468852 687254
rect 468568 687012 468622 687176
rect 468622 687012 468806 687176
rect 468806 687012 468852 687176
rect 468568 686950 468852 687012
rect 512924 686746 517294 691578
rect 519782 686746 524152 691578
rect 222764 656624 224356 664238
rect 442366 656090 442650 656156
rect 442366 655926 442412 656090
rect 442412 655926 442596 656090
rect 442596 655926 442650 656090
rect 442366 655852 442650 655926
rect 442760 656090 443044 656164
rect 442760 655926 442812 656090
rect 442812 655926 442996 656090
rect 442996 655926 443044 656090
rect 442760 655860 443044 655926
rect 442356 655290 442684 655372
rect 442356 655126 442412 655290
rect 442412 655126 442596 655290
rect 442596 655126 442684 655290
rect 442356 655076 442684 655126
rect 442768 655290 443052 655368
rect 442768 655126 442822 655290
rect 442822 655126 443006 655290
rect 443006 655126 443052 655290
rect 442768 655064 443052 655126
rect 450766 656090 451050 656156
rect 450766 655926 450812 656090
rect 450812 655926 450996 656090
rect 450996 655926 451050 656090
rect 450766 655852 451050 655926
rect 451160 656090 451444 656164
rect 451160 655926 451212 656090
rect 451212 655926 451396 656090
rect 451396 655926 451444 656090
rect 451160 655860 451444 655926
rect 450756 655290 451084 655372
rect 450756 655126 450812 655290
rect 450812 655126 450996 655290
rect 450996 655126 451084 655290
rect 450756 655076 451084 655126
rect 451168 655290 451452 655368
rect 451168 655126 451222 655290
rect 451222 655126 451406 655290
rect 451406 655126 451452 655290
rect 451168 655064 451452 655126
rect 134622 596998 135400 597544
rect 135822 596998 136600 597544
rect 137022 596998 137800 597544
rect 138222 596998 139000 597544
rect 85622 582998 86400 583544
rect 86822 582998 87600 583544
rect 88022 582998 88800 583544
rect 89222 582998 90000 583544
rect 416472 586394 417092 586782
rect 416472 584684 417092 585072
rect 101632 565036 102410 565582
rect 102832 565036 103610 565582
rect 104032 565036 104810 565582
rect 105232 565036 106010 565582
rect 107622 564998 108400 565544
rect 108822 564998 109600 565544
rect 110022 564998 110800 565544
rect 111222 564998 112000 565544
<< metal5 >>
rect 165594 702540 170594 704800
rect 165552 702300 170594 702540
rect 175894 702434 180894 704800
rect 175862 702300 180894 702434
rect 217294 702970 222294 704800
rect 217294 702300 222336 702970
rect 227594 702926 232594 704800
rect 31620 696030 43302 698312
rect 165552 696162 170568 702300
rect 31620 695992 112194 696030
rect 31620 695542 118390 695992
rect 31620 694458 116918 695542
rect 118020 694458 118390 695542
rect 31620 694138 118390 694458
rect 31620 694130 112194 694138
rect 31620 680316 43302 694130
rect 165552 693934 170584 696162
rect 165554 682686 170584 693934
rect 175862 682686 180868 702300
rect 217306 684124 222336 702300
rect 165508 682660 187874 682686
rect 217280 682660 222336 684124
rect 227582 694624 232594 702926
rect 318994 702300 323994 704800
rect 329294 702300 334294 704800
rect 227582 682660 232548 694624
rect 511622 691578 524830 694392
rect 416118 688050 416878 688698
rect 416118 688042 416560 688050
rect 416118 687738 416166 688042
rect 416450 687746 416560 688042
rect 416844 687850 416878 688050
rect 468118 688052 468878 688698
rect 473182 688052 474038 688056
rect 468118 688050 474038 688052
rect 468118 688042 468560 688050
rect 416844 687746 420894 687850
rect 416450 687738 420894 687746
rect 416118 687298 420894 687738
rect 416118 687258 416878 687298
rect 416118 686962 416156 687258
rect 416484 687254 416878 687258
rect 416484 686962 416568 687254
rect 416118 686950 416568 686962
rect 416852 686950 416878 687254
rect 416118 686838 416878 686950
rect 420072 686994 420894 687298
rect 468118 687738 468166 688042
rect 468450 687746 468560 688042
rect 468844 687746 474038 688050
rect 468450 687738 474038 687746
rect 468118 687500 474038 687738
rect 468118 687298 468896 687500
rect 468118 687258 468878 687298
rect 420072 685576 420916 686994
rect 468118 686962 468156 687258
rect 468484 687254 468878 687258
rect 468484 686962 468568 687254
rect 468118 686950 468568 686962
rect 468852 686950 468878 687254
rect 468118 686838 468878 686950
rect 473182 686592 474038 687500
rect 511622 686746 512924 691578
rect 517294 686746 519782 691578
rect 524152 686746 524830 691578
rect 165508 682658 191410 682660
rect 208250 682658 232548 682660
rect 31582 663992 43430 680316
rect 165508 677212 191570 682658
rect 185918 677168 191570 677212
rect 31582 663542 66390 663992
rect 31582 662458 64918 663542
rect 66020 662458 66390 663542
rect 31582 662138 66390 662458
rect 31582 552010 43430 662138
rect 134234 597778 139152 597946
rect 134182 597544 139154 597778
rect 134182 596998 134622 597544
rect 135400 596998 135822 597544
rect 136600 596998 137022 597544
rect 137800 596998 138222 597544
rect 139000 596998 139154 597544
rect 134182 596126 139154 596998
rect 134182 595332 139146 596126
rect 134076 592180 139146 595332
rect 85234 583778 90152 583946
rect 85182 583544 90154 583778
rect 85182 582998 85622 583544
rect 86400 582998 86822 583544
rect 87600 582998 88022 583544
rect 88800 582998 89222 583544
rect 90000 582998 90154 583544
rect 85182 580040 90154 582998
rect 85182 576158 90162 580040
rect 85182 569934 90170 576158
rect 85182 552010 90102 569934
rect 101244 565954 106156 565984
rect 101244 565946 108222 565954
rect 101244 565816 112152 565946
rect 101238 565778 112152 565816
rect 101238 565582 112154 565778
rect 101238 565036 101632 565582
rect 102410 565036 102832 565582
rect 103610 565036 104032 565582
rect 104810 565036 105232 565582
rect 106010 565544 112154 565582
rect 106010 565036 107622 565544
rect 101238 564998 107622 565036
rect 108400 564998 108822 565544
rect 109600 564998 110022 565544
rect 110800 564998 111222 565544
rect 112000 564998 112154 565544
rect 101238 564532 112154 564998
rect 101184 564454 112154 564532
rect 31582 551954 93230 552010
rect 101184 551954 112166 564454
rect 134076 551954 139428 592180
rect 186722 585092 191570 677168
rect 204138 677168 232548 682658
rect 420086 681318 420914 685576
rect 265894 681262 420914 681318
rect 247820 681228 420914 681262
rect 473190 681228 474018 686592
rect 511622 681228 524830 686746
rect 247820 677672 524916 681228
rect 247820 677366 420902 677672
rect 247820 677310 275360 677366
rect 204138 591614 209704 677168
rect 222390 664238 224726 664668
rect 222390 656624 222764 664238
rect 224356 662136 224726 664238
rect 247820 662136 252154 677310
rect 224356 658694 252154 662136
rect 224356 656624 224726 658694
rect 247820 658682 252154 658694
rect 444102 656820 444930 677672
rect 453478 656822 454306 677672
rect 452080 656820 454306 656822
rect 222390 656366 224726 656624
rect 442316 656164 444930 656820
rect 442316 656156 442760 656164
rect 442316 655852 442366 656156
rect 442650 655860 442760 656156
rect 443044 655860 444930 656164
rect 442650 655852 444930 655860
rect 442316 655372 444930 655852
rect 442316 655076 442356 655372
rect 442684 655368 444930 655372
rect 442684 655076 442768 655368
rect 442316 655064 442768 655076
rect 443052 655064 444930 655368
rect 442316 654954 444930 655064
rect 450716 656164 454306 656820
rect 450716 656156 451160 656164
rect 450716 655852 450766 656156
rect 451050 655860 451160 656156
rect 451444 655860 454306 656164
rect 451050 655852 454306 655860
rect 450716 655372 454306 655852
rect 450716 655076 450756 655372
rect 451084 655368 454306 655372
rect 451084 655076 451168 655368
rect 450716 655064 451168 655076
rect 451452 655064 454306 655368
rect 450716 654954 454306 655064
rect 442318 654952 443078 654954
rect 444102 650610 444930 654954
rect 450718 654952 451478 654954
rect 452080 654944 454306 654954
rect 453478 650320 454306 654944
rect 204098 590968 209704 591614
rect 204098 588300 209692 590968
rect 204114 587926 209692 588300
rect 204114 587886 211476 587926
rect 402686 587900 410794 587910
rect 414686 587900 417000 587904
rect 402686 587886 417000 587900
rect 204114 587862 218504 587886
rect 230148 587862 417000 587886
rect 204114 587396 417000 587862
rect 204114 587374 233540 587396
rect 402686 587378 417000 587396
rect 204114 587372 211476 587374
rect 204114 586508 209692 587372
rect 410316 587368 417000 587378
rect 416544 587070 417000 587368
rect 416544 586912 417002 587070
rect 416354 586782 417192 586912
rect 416354 586394 416472 586782
rect 417092 586394 417192 586782
rect 416354 586296 417192 586394
rect 186716 584756 191570 585092
rect 416354 585072 417186 585172
rect 186716 583460 191564 584756
rect 416354 584684 416472 585072
rect 417092 584684 417186 585072
rect 416354 584586 417186 584684
rect 416574 583490 416992 584586
rect 410490 583488 416992 583490
rect 404554 583468 416992 583488
rect 223084 583460 416992 583468
rect 186716 582996 416992 583460
rect 223084 582978 416992 582996
rect 404554 582974 416836 582978
rect 404554 582972 410596 582974
rect 417360 582210 424026 583390
rect 417360 582198 423992 582210
rect 417360 581742 423936 582198
rect 417360 581570 424026 581742
rect 417350 580238 424026 581570
rect 417358 579200 424026 580238
rect 417358 551998 423994 579200
rect 511622 554468 524830 677672
rect 511624 552106 524830 554468
rect 417276 551954 476240 551998
rect 31582 551888 476240 551954
rect 511624 551896 524886 552106
rect 499162 551888 524886 551896
rect 31582 542478 524886 551888
rect 31582 542438 433714 542478
rect 499162 542446 524886 542478
rect 31656 542384 433714 542438
rect 31656 542284 93230 542384
<< comment >>
rect -100 704000 584100 704100
rect -100 0 0 704000
rect 584000 0 584100 704000
rect -100 -100 584100 0
use comparator_v6  comparator_v6_0
timestamp 1654337383
transform 0 1 419266 1 0 584802
box -2598 -1934 4390 5556
use sky130_fd_pr__diode_pd2nw_05v5_RT56W3  sky130_fd_pr__diode_pd2nw_05v5_RT56W3_0
timestamp 1654421061
transform 1 0 74128 0 1 662860
box -321 -321 321 321
use sky130_fd_pr__diode_pd2nw_05v5_RT56W3  sky130_fd_pr__diode_pd2nw_05v5_RT56W3_1
timestamp 1654421061
transform 1 0 126100 0 1 694854
box -321 -321 321 321
use sky130_fd_pr__diode_pw2nd_05v5_GT7E3L  sky130_fd_pr__diode_pw2nd_05v5_GT7E3L_0
timestamp 1654419227
transform 1 0 67028 0 1 663058
box -183 -183 183 183
use sky130_fd_pr__diode_pw2nd_05v5_GT7G3L  sky130_fd_pr__diode_pw2nd_05v5_GT7G3L_0
timestamp 1654421061
transform 1 0 118990 0 1 695058
box -183 -183 183 183
use sky130_fd_sc_hd__buf_2  sky130_fd_sc_hd__buf_2_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1654337383
transform 1 0 85632 0 1 585240
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  sky130_fd_sc_hd__buf_2_1
timestamp 1654337383
transform 1 0 103250 0 1 567442
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  sky130_fd_sc_hd__buf_2_2
timestamp 1654337383
transform 1 0 134624 0 1 599244
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  sky130_fd_sc_hd__buf_2_3
timestamp 1654337383
transform 0 -1 440656 1 0 655486
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  sky130_fd_sc_hd__buf_2_4
timestamp 1654337383
transform 0 -1 449242 1 0 655494
box -38 -48 406 592
use sky130_fd_sc_hd__buf_16  sky130_fd_sc_hd__buf_16_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1654337383
transform 1 0 87054 0 1 585244
box -38 -48 2062 592
use sky130_fd_sc_hd__buf_16  sky130_fd_sc_hd__buf_16_1
timestamp 1654337383
transform 1 0 108006 0 1 567526
box -38 -48 2062 592
use sky130_fd_sc_hd__buf_16  sky130_fd_sc_hd__buf_16_2
timestamp 1654337383
transform 1 0 136168 0 1 599250
box -38 -48 2062 592
use sky130_fd_sc_hd__buf_16  sky130_fd_sc_hd__buf_16_3
timestamp 1654337383
transform 0 -1 415762 1 0 686886
box -38 -48 2062 592
use sky130_fd_sc_hd__buf_16  sky130_fd_sc_hd__buf_16_4
timestamp 1654337383
transform 0 -1 467696 1 0 686840
box -38 -48 2062 592
<< labels >>
flabel metal3 s 583520 269230 584800 269342 0 FreeSans 1120 0 0 0 gpio_analog[0]
port 0 nsew signal bidirectional
flabel metal3 s -800 381864 480 381976 0 FreeSans 1120 0 0 0 gpio_analog[10]
port 1 nsew signal bidirectional
flabel metal3 s -800 338642 480 338754 0 FreeSans 1120 0 0 0 gpio_analog[11]
port 2 nsew signal bidirectional
flabel metal3 s -800 295420 480 295532 0 FreeSans 1120 0 0 0 gpio_analog[12]
port 3 nsew signal bidirectional
flabel metal3 s -800 252398 480 252510 0 FreeSans 1120 0 0 0 gpio_analog[13]
port 4 nsew signal bidirectional
flabel metal3 s -800 124776 480 124888 0 FreeSans 1120 0 0 0 gpio_analog[14]
port 5 nsew signal bidirectional
flabel metal3 s -800 81554 480 81666 0 FreeSans 1120 0 0 0 gpio_analog[15]
port 6 nsew signal bidirectional
flabel metal3 s -800 38332 480 38444 0 FreeSans 1120 0 0 0 gpio_analog[16]
port 7 nsew signal bidirectional
flabel metal3 s -800 16910 480 17022 0 FreeSans 1120 0 0 0 gpio_analog[17]
port 8 nsew signal bidirectional
flabel metal3 s 583520 313652 584800 313764 0 FreeSans 1120 0 0 0 gpio_analog[1]
port 9 nsew signal bidirectional
flabel metal3 s 583520 358874 584800 358986 0 FreeSans 1120 0 0 0 gpio_analog[2]
port 10 nsew signal bidirectional
flabel metal3 s 583520 405296 584800 405408 0 FreeSans 1120 0 0 0 gpio_analog[3]
port 11 nsew signal bidirectional
flabel metal3 s 583520 449718 584800 449830 0 FreeSans 1120 0 0 0 gpio_analog[4]
port 12 nsew signal bidirectional
flabel metal3 s 583520 494140 584800 494252 0 FreeSans 1120 0 0 0 gpio_analog[5]
port 13 nsew signal bidirectional
flabel metal3 s 583520 583562 584800 583674 0 FreeSans 1120 0 0 0 gpio_analog[6]
port 14 nsew signal bidirectional
flabel metal3 s -800 511530 480 511642 0 FreeSans 1120 0 0 0 gpio_analog[7]
port 15 nsew signal bidirectional
flabel metal3 s -800 468308 480 468420 0 FreeSans 1120 0 0 0 gpio_analog[8]
port 16 nsew signal bidirectional
flabel metal3 s -800 425086 480 425198 0 FreeSans 1120 0 0 0 gpio_analog[9]
port 17 nsew signal bidirectional
flabel metal3 s 583520 270412 584800 270524 0 FreeSans 1120 0 0 0 gpio_noesd[0]
port 18 nsew signal bidirectional
flabel metal3 s -800 380682 480 380794 0 FreeSans 1120 0 0 0 gpio_noesd[10]
port 19 nsew signal bidirectional
flabel metal3 s -800 337460 480 337572 0 FreeSans 1120 0 0 0 gpio_noesd[11]
port 20 nsew signal bidirectional
flabel metal3 s -800 294238 480 294350 0 FreeSans 1120 0 0 0 gpio_noesd[12]
port 21 nsew signal bidirectional
flabel metal3 s -800 251216 480 251328 0 FreeSans 1120 0 0 0 gpio_noesd[13]
port 22 nsew signal bidirectional
flabel metal3 s -800 123594 480 123706 0 FreeSans 1120 0 0 0 gpio_noesd[14]
port 23 nsew signal bidirectional
flabel metal3 s -800 80372 480 80484 0 FreeSans 1120 0 0 0 gpio_noesd[15]
port 24 nsew signal bidirectional
flabel metal3 s -800 37150 480 37262 0 FreeSans 1120 0 0 0 gpio_noesd[16]
port 25 nsew signal bidirectional
flabel metal3 s -800 15728 480 15840 0 FreeSans 1120 0 0 0 gpio_noesd[17]
port 26 nsew signal bidirectional
flabel metal3 s 583520 314834 584800 314946 0 FreeSans 1120 0 0 0 gpio_noesd[1]
port 27 nsew signal bidirectional
flabel metal3 s 583520 360056 584800 360168 0 FreeSans 1120 0 0 0 gpio_noesd[2]
port 28 nsew signal bidirectional
flabel metal3 s 583520 406478 584800 406590 0 FreeSans 1120 0 0 0 gpio_noesd[3]
port 29 nsew signal bidirectional
flabel metal3 s 583520 450900 584800 451012 0 FreeSans 1120 0 0 0 gpio_noesd[4]
port 30 nsew signal bidirectional
flabel metal3 s 583520 495322 584800 495434 0 FreeSans 1120 0 0 0 gpio_noesd[5]
port 31 nsew signal bidirectional
flabel metal3 s 583520 584744 584800 584856 0 FreeSans 1120 0 0 0 gpio_noesd[6]
port 32 nsew signal bidirectional
flabel metal3 s -800 510348 480 510460 0 FreeSans 1120 0 0 0 gpio_noesd[7]
port 33 nsew signal bidirectional
flabel metal3 s -800 467126 480 467238 0 FreeSans 1120 0 0 0 gpio_noesd[8]
port 34 nsew signal bidirectional
flabel metal3 s -800 423904 480 424016 0 FreeSans 1120 0 0 0 gpio_noesd[9]
port 35 nsew signal bidirectional
flabel metal3 s 582300 677984 584800 682984 0 FreeSans 1120 0 0 0 io_analog[0]
port 36 nsew signal bidirectional
flabel metal3 s 0 680242 1700 685242 0 FreeSans 1120 0 0 0 io_analog[10]
port 37 nsew signal bidirectional
flabel metal3 s 566594 702300 571594 704800 0 FreeSans 1920 180 0 0 io_analog[1]
port 38 nsew signal bidirectional
flabel metal3 s 465394 702300 470394 704800 0 FreeSans 1920 180 0 0 io_analog[2]
port 39 nsew signal bidirectional
flabel metal3 s 413394 702300 418394 704800 0 FreeSans 1920 180 0 0 io_analog[3]
port 40 nsew signal bidirectional
flabel metal3 s 329294 702300 334294 704800 0 FreeSans 1920 180 0 0 io_analog[4]
port 41 nsew signal bidirectional
flabel metal4 s 329294 702300 334294 704800 0 FreeSans 1920 180 0 0 io_analog[4]
port 41 nsew signal bidirectional
flabel metal5 s 329294 702300 334294 704800 0 FreeSans 1920 180 0 0 io_analog[4]
port 41 nsew signal bidirectional
flabel metal3 s 227594 702300 232594 704800 0 FreeSans 1920 180 0 0 io_analog[5]
port 42 nsew signal bidirectional
flabel metal4 s 227594 702300 232594 704800 0 FreeSans 1920 180 0 0 io_analog[5]
port 42 nsew signal bidirectional
flabel metal5 s 227594 702300 232594 704800 0 FreeSans 1920 180 0 0 io_analog[5]
port 42 nsew signal bidirectional
flabel metal3 s 175894 702300 180894 704800 0 FreeSans 1920 180 0 0 io_analog[6]
port 43 nsew signal bidirectional
flabel metal4 s 175894 702300 180894 704800 0 FreeSans 1920 180 0 0 io_analog[6]
port 43 nsew signal bidirectional
flabel metal5 s 175894 702300 180894 704800 0 FreeSans 1920 180 0 0 io_analog[6]
port 43 nsew signal bidirectional
flabel metal3 s 68194 702300 73194 704800 0 FreeSans 1920 180 0 0 io_analog[8]
port 45 nsew signal bidirectional
flabel metal3 s 16194 702300 21194 704800 0 FreeSans 1920 180 0 0 io_analog[9]
port 46 nsew signal bidirectional
flabel metal3 s 318994 702300 323994 704800 0 FreeSans 1920 180 0 0 io_analog[4]
port 47 nsew signal bidirectional
flabel metal4 s 318994 702300 323994 704800 0 FreeSans 1920 180 0 0 io_analog[4]
port 47 nsew signal bidirectional
flabel metal5 s 318994 702300 323994 704800 0 FreeSans 1920 180 0 0 io_analog[4]
port 47 nsew signal bidirectional
flabel metal3 s 217294 702300 222294 704800 0 FreeSans 1920 180 0 0 io_analog[5]
port 48 nsew signal bidirectional
flabel metal4 s 217294 702300 222294 704800 0 FreeSans 1920 180 0 0 io_analog[5]
port 48 nsew signal bidirectional
flabel metal5 s 217294 702300 222294 704800 0 FreeSans 1920 180 0 0 io_analog[5]
port 48 nsew signal bidirectional
flabel metal3 s 165594 702300 170594 704800 0 FreeSans 1920 180 0 0 io_analog[6]
port 49 nsew signal bidirectional
flabel metal4 s 165594 702300 170594 704800 0 FreeSans 1920 180 0 0 io_analog[6]
port 49 nsew signal bidirectional
flabel metal5 s 165594 702300 170594 704800 0 FreeSans 1920 180 0 0 io_analog[6]
port 49 nsew signal bidirectional
flabel metal3 s 326794 702300 328994 704800 0 FreeSans 1920 180 0 0 io_clamp_high[0]
port 50 nsew signal bidirectional
flabel metal3 s 225094 702300 227294 704800 0 FreeSans 1920 180 0 0 io_clamp_high[1]
port 51 nsew signal bidirectional
flabel metal3 s 173394 702300 175594 704800 0 FreeSans 1920 180 0 0 io_clamp_high[2]
port 52 nsew signal bidirectional
flabel metal3 s 324294 702300 326494 704800 0 FreeSans 1920 180 0 0 io_clamp_low[0]
port 53 nsew signal bidirectional
flabel metal3 s 222594 702300 224794 704800 0 FreeSans 1920 180 0 0 io_clamp_low[1]
port 54 nsew signal bidirectional
flabel metal3 s 170894 702300 173094 704800 0 FreeSans 1920 180 0 0 io_clamp_low[2]
port 55 nsew signal bidirectional
flabel metal3 s 583520 2726 584800 2838 0 FreeSans 1120 0 0 0 io_in[0]
port 56 nsew signal input
flabel metal3 s 583520 408842 584800 408954 0 FreeSans 1120 0 0 0 io_in[10]
port 57 nsew signal input
flabel metal3 s 583520 453264 584800 453376 0 FreeSans 1120 0 0 0 io_in[11]
port 58 nsew signal input
flabel metal3 s 583520 497686 584800 497798 0 FreeSans 1120 0 0 0 io_in[12]
port 59 nsew signal input
flabel metal3 s 583520 587108 584800 587220 0 FreeSans 1120 0 0 0 io_in[13]
port 60 nsew signal input
flabel metal3 s -800 507984 480 508096 0 FreeSans 1120 0 0 0 io_in[14]
port 61 nsew signal input
flabel metal3 s -800 464762 480 464874 0 FreeSans 1120 0 0 0 io_in[15]
port 62 nsew signal input
flabel metal3 s -800 421540 480 421652 0 FreeSans 1120 0 0 0 io_in[16]
port 63 nsew signal input
flabel metal3 s -800 378318 480 378430 0 FreeSans 1120 0 0 0 io_in[17]
port 64 nsew signal input
flabel metal3 s -800 335096 480 335208 0 FreeSans 1120 0 0 0 io_in[18]
port 65 nsew signal input
flabel metal3 s -800 291874 480 291986 0 FreeSans 1120 0 0 0 io_in[19]
port 66 nsew signal input
flabel metal3 s 583520 7454 584800 7566 0 FreeSans 1120 0 0 0 io_in[1]
port 67 nsew signal input
flabel metal3 s -800 248852 480 248964 0 FreeSans 1120 0 0 0 io_in[20]
port 68 nsew signal input
flabel metal3 s -800 121230 480 121342 0 FreeSans 1120 0 0 0 io_in[21]
port 69 nsew signal input
flabel metal3 s -800 78008 480 78120 0 FreeSans 1120 0 0 0 io_in[22]
port 70 nsew signal input
flabel metal3 s -800 34786 480 34898 0 FreeSans 1120 0 0 0 io_in[23]
port 71 nsew signal input
flabel metal3 s -800 13364 480 13476 0 FreeSans 1120 0 0 0 io_in[24]
port 72 nsew signal input
flabel metal3 s -800 8636 480 8748 0 FreeSans 1120 0 0 0 io_in[25]
port 73 nsew signal input
flabel metal3 s -800 3908 480 4020 0 FreeSans 1120 0 0 0 io_in[26]
port 74 nsew signal input
flabel metal3 s 583520 12182 584800 12294 0 FreeSans 1120 0 0 0 io_in[2]
port 75 nsew signal input
flabel metal3 s 583520 16910 584800 17022 0 FreeSans 1120 0 0 0 io_in[3]
port 76 nsew signal input
flabel metal3 s 583520 21638 584800 21750 0 FreeSans 1120 0 0 0 io_in[4]
port 77 nsew signal input
flabel metal3 s 583520 48096 584800 48208 0 FreeSans 1120 0 0 0 io_in[5]
port 78 nsew signal input
flabel metal3 s 583520 92754 584800 92866 0 FreeSans 1120 0 0 0 io_in[6]
port 79 nsew signal input
flabel metal3 s 583520 272776 584800 272888 0 FreeSans 1120 0 0 0 io_in[7]
port 80 nsew signal input
flabel metal3 s 583520 317198 584800 317310 0 FreeSans 1120 0 0 0 io_in[8]
port 81 nsew signal input
flabel metal3 s 583520 362420 584800 362532 0 FreeSans 1120 0 0 0 io_in[9]
port 82 nsew signal input
flabel metal3 s 583520 1544 584800 1656 0 FreeSans 1120 0 0 0 io_in_3v3[0]
port 83 nsew signal input
flabel metal3 s 583520 407660 584800 407772 0 FreeSans 1120 0 0 0 io_in_3v3[10]
port 84 nsew signal input
flabel metal3 s 583520 452082 584800 452194 0 FreeSans 1120 0 0 0 io_in_3v3[11]
port 85 nsew signal input
flabel metal3 s 583520 496504 584800 496616 0 FreeSans 1120 0 0 0 io_in_3v3[12]
port 86 nsew signal input
flabel metal3 s 583520 585926 584800 586038 0 FreeSans 1120 0 0 0 io_in_3v3[13]
port 87 nsew signal input
flabel metal3 s -800 509166 480 509278 0 FreeSans 1120 0 0 0 io_in_3v3[14]
port 88 nsew signal input
flabel metal3 s -800 465944 480 466056 0 FreeSans 1120 0 0 0 io_in_3v3[15]
port 89 nsew signal input
flabel metal3 s -800 422722 480 422834 0 FreeSans 1120 0 0 0 io_in_3v3[16]
port 90 nsew signal input
flabel metal3 s -800 379500 480 379612 0 FreeSans 1120 0 0 0 io_in_3v3[17]
port 91 nsew signal input
flabel metal3 s -800 336278 480 336390 0 FreeSans 1120 0 0 0 io_in_3v3[18]
port 92 nsew signal input
flabel metal3 s -800 293056 480 293168 0 FreeSans 1120 0 0 0 io_in_3v3[19]
port 93 nsew signal input
flabel metal3 s 583520 6272 584800 6384 0 FreeSans 1120 0 0 0 io_in_3v3[1]
port 94 nsew signal input
flabel metal3 s -800 250034 480 250146 0 FreeSans 1120 0 0 0 io_in_3v3[20]
port 95 nsew signal input
flabel metal3 s -800 122412 480 122524 0 FreeSans 1120 0 0 0 io_in_3v3[21]
port 96 nsew signal input
flabel metal3 s -800 79190 480 79302 0 FreeSans 1120 0 0 0 io_in_3v3[22]
port 97 nsew signal input
flabel metal3 s -800 35968 480 36080 0 FreeSans 1120 0 0 0 io_in_3v3[23]
port 98 nsew signal input
flabel metal3 s -800 14546 480 14658 0 FreeSans 1120 0 0 0 io_in_3v3[24]
port 99 nsew signal input
flabel metal3 s -800 9818 480 9930 0 FreeSans 1120 0 0 0 io_in_3v3[25]
port 100 nsew signal input
flabel metal3 s -800 5090 480 5202 0 FreeSans 1120 0 0 0 io_in_3v3[26]
port 101 nsew signal input
flabel metal3 s 583520 11000 584800 11112 0 FreeSans 1120 0 0 0 io_in_3v3[2]
port 102 nsew signal input
flabel metal3 s 583520 15728 584800 15840 0 FreeSans 1120 0 0 0 io_in_3v3[3]
port 103 nsew signal input
flabel metal3 s 583520 20456 584800 20568 0 FreeSans 1120 0 0 0 io_in_3v3[4]
port 104 nsew signal input
flabel metal3 s 583520 46914 584800 47026 0 FreeSans 1120 0 0 0 io_in_3v3[5]
port 105 nsew signal input
flabel metal3 s 583520 91572 584800 91684 0 FreeSans 1120 0 0 0 io_in_3v3[6]
port 106 nsew signal input
flabel metal3 s 583520 271594 584800 271706 0 FreeSans 1120 0 0 0 io_in_3v3[7]
port 107 nsew signal input
flabel metal3 s 583520 316016 584800 316128 0 FreeSans 1120 0 0 0 io_in_3v3[8]
port 108 nsew signal input
flabel metal3 s 583520 361238 584800 361350 0 FreeSans 1120 0 0 0 io_in_3v3[9]
port 109 nsew signal input
flabel metal3 s 583520 5090 584800 5202 0 FreeSans 1120 0 0 0 io_oeb[0]
port 110 nsew signal tristate
flabel metal3 s 583520 411206 584800 411318 0 FreeSans 1120 0 0 0 io_oeb[10]
port 111 nsew signal tristate
flabel metal3 s 583520 455628 584800 455740 0 FreeSans 1120 0 0 0 io_oeb[11]
port 112 nsew signal tristate
flabel metal3 s 583520 500050 584800 500162 0 FreeSans 1120 0 0 0 io_oeb[12]
port 113 nsew signal tristate
flabel metal3 s 583520 589472 584800 589584 0 FreeSans 1120 0 0 0 io_oeb[13]
port 114 nsew signal tristate
flabel metal3 s -800 505620 480 505732 0 FreeSans 1120 0 0 0 io_oeb[14]
port 115 nsew signal tristate
flabel metal3 s -800 462398 480 462510 0 FreeSans 1120 0 0 0 io_oeb[15]
port 116 nsew signal tristate
flabel metal3 s -800 419176 480 419288 0 FreeSans 1120 0 0 0 io_oeb[16]
port 117 nsew signal tristate
flabel metal3 s -800 375954 480 376066 0 FreeSans 1120 0 0 0 io_oeb[17]
port 118 nsew signal tristate
flabel metal3 s -800 332732 480 332844 0 FreeSans 1120 0 0 0 io_oeb[18]
port 119 nsew signal tristate
flabel metal3 s -800 289510 480 289622 0 FreeSans 1120 0 0 0 io_oeb[19]
port 120 nsew signal tristate
flabel metal3 s 583520 9818 584800 9930 0 FreeSans 1120 0 0 0 io_oeb[1]
port 121 nsew signal tristate
flabel metal3 s -800 246488 480 246600 0 FreeSans 1120 0 0 0 io_oeb[20]
port 122 nsew signal tristate
flabel metal3 s -800 118866 480 118978 0 FreeSans 1120 0 0 0 io_oeb[21]
port 123 nsew signal tristate
flabel metal3 s -800 75644 480 75756 0 FreeSans 1120 0 0 0 io_oeb[22]
port 124 nsew signal tristate
flabel metal3 s -800 32422 480 32534 0 FreeSans 1120 0 0 0 io_oeb[23]
port 125 nsew signal tristate
flabel metal3 s -800 11000 480 11112 0 FreeSans 1120 0 0 0 io_oeb[24]
port 126 nsew signal tristate
flabel metal3 s -800 6272 480 6384 0 FreeSans 1120 0 0 0 io_oeb[25]
port 127 nsew signal tristate
flabel metal3 s -800 1544 480 1656 0 FreeSans 1120 0 0 0 io_oeb[26]
port 128 nsew signal tristate
flabel metal3 s 583520 14546 584800 14658 0 FreeSans 1120 0 0 0 io_oeb[2]
port 129 nsew signal tristate
flabel metal3 s 583520 19274 584800 19386 0 FreeSans 1120 0 0 0 io_oeb[3]
port 130 nsew signal tristate
flabel metal3 s 583520 24002 584800 24114 0 FreeSans 1120 0 0 0 io_oeb[4]
port 131 nsew signal tristate
flabel metal3 s 583520 50460 584800 50572 0 FreeSans 1120 0 0 0 io_oeb[5]
port 132 nsew signal tristate
flabel metal3 s 583520 95118 584800 95230 0 FreeSans 1120 0 0 0 io_oeb[6]
port 133 nsew signal tristate
flabel metal3 s 583520 275140 584800 275252 0 FreeSans 1120 0 0 0 io_oeb[7]
port 134 nsew signal tristate
flabel metal3 s 583520 319562 584800 319674 0 FreeSans 1120 0 0 0 io_oeb[8]
port 135 nsew signal tristate
flabel metal3 s 583520 364784 584800 364896 0 FreeSans 1120 0 0 0 io_oeb[9]
port 136 nsew signal tristate
flabel metal3 s 583520 3908 584800 4020 0 FreeSans 1120 0 0 0 io_out[0]
port 137 nsew signal tristate
flabel metal3 s 583520 410024 584800 410136 0 FreeSans 1120 0 0 0 io_out[10]
port 138 nsew signal tristate
flabel metal3 s 583520 454446 584800 454558 0 FreeSans 1120 0 0 0 io_out[11]
port 139 nsew signal tristate
flabel metal3 s 583520 498868 584800 498980 0 FreeSans 1120 0 0 0 io_out[12]
port 140 nsew signal tristate
flabel metal3 s 583520 588290 584800 588402 0 FreeSans 1120 0 0 0 io_out[13]
port 141 nsew signal tristate
flabel metal3 s -800 506802 480 506914 0 FreeSans 1120 0 0 0 io_out[14]
port 142 nsew signal tristate
flabel metal3 s -800 463580 480 463692 0 FreeSans 1120 0 0 0 io_out[15]
port 143 nsew signal tristate
flabel metal3 s -800 420358 480 420470 0 FreeSans 1120 0 0 0 io_out[16]
port 144 nsew signal tristate
flabel metal3 s -800 377136 480 377248 0 FreeSans 1120 0 0 0 io_out[17]
port 145 nsew signal tristate
flabel metal3 s -800 333914 480 334026 0 FreeSans 1120 0 0 0 io_out[18]
port 146 nsew signal tristate
flabel metal3 s -800 290692 480 290804 0 FreeSans 1120 0 0 0 io_out[19]
port 147 nsew signal tristate
flabel metal3 s 583520 8636 584800 8748 0 FreeSans 1120 0 0 0 io_out[1]
port 148 nsew signal tristate
flabel metal3 s -800 247670 480 247782 0 FreeSans 1120 0 0 0 io_out[20]
port 149 nsew signal tristate
flabel metal3 s -800 120048 480 120160 0 FreeSans 1120 0 0 0 io_out[21]
port 150 nsew signal tristate
flabel metal3 s -800 76826 480 76938 0 FreeSans 1120 0 0 0 io_out[22]
port 151 nsew signal tristate
flabel metal3 s -800 33604 480 33716 0 FreeSans 1120 0 0 0 io_out[23]
port 152 nsew signal tristate
flabel metal3 s -800 12182 480 12294 0 FreeSans 1120 0 0 0 io_out[24]
port 153 nsew signal tristate
flabel metal3 s -800 7454 480 7566 0 FreeSans 1120 0 0 0 io_out[25]
port 154 nsew signal tristate
flabel metal3 s -800 2726 480 2838 0 FreeSans 1120 0 0 0 io_out[26]
port 155 nsew signal tristate
flabel metal3 s 583520 13364 584800 13476 0 FreeSans 1120 0 0 0 io_out[2]
port 156 nsew signal tristate
flabel metal3 s 583520 18092 584800 18204 0 FreeSans 1120 0 0 0 io_out[3]
port 157 nsew signal tristate
flabel metal3 s 583520 22820 584800 22932 0 FreeSans 1120 0 0 0 io_out[4]
port 158 nsew signal tristate
flabel metal3 s 583520 49278 584800 49390 0 FreeSans 1120 0 0 0 io_out[5]
port 159 nsew signal tristate
flabel metal3 s 583520 93936 584800 94048 0 FreeSans 1120 0 0 0 io_out[6]
port 160 nsew signal tristate
flabel metal3 s 583520 273958 584800 274070 0 FreeSans 1120 0 0 0 io_out[7]
port 161 nsew signal tristate
flabel metal3 s 583520 318380 584800 318492 0 FreeSans 1120 0 0 0 io_out[8]
port 162 nsew signal tristate
flabel metal3 s 583520 363602 584800 363714 0 FreeSans 1120 0 0 0 io_out[9]
port 163 nsew signal tristate
flabel metal2 s 125816 -800 125928 480 0 FreeSans 1120 90 0 0 la_data_in[0]
port 164 nsew signal input
flabel metal2 s 480416 -800 480528 480 0 FreeSans 1120 90 0 0 la_data_in[100]
port 165 nsew signal input
flabel metal2 s 483962 -800 484074 480 0 FreeSans 1120 90 0 0 la_data_in[101]
port 166 nsew signal input
flabel metal2 s 487508 -800 487620 480 0 FreeSans 1120 90 0 0 la_data_in[102]
port 167 nsew signal input
flabel metal2 s 491054 -800 491166 480 0 FreeSans 1120 90 0 0 la_data_in[103]
port 168 nsew signal input
flabel metal2 s 494600 -800 494712 480 0 FreeSans 1120 90 0 0 la_data_in[104]
port 169 nsew signal input
flabel metal2 s 498146 -800 498258 480 0 FreeSans 1120 90 0 0 la_data_in[105]
port 170 nsew signal input
flabel metal2 s 501692 -800 501804 480 0 FreeSans 1120 90 0 0 la_data_in[106]
port 171 nsew signal input
flabel metal2 s 505238 -800 505350 480 0 FreeSans 1120 90 0 0 la_data_in[107]
port 172 nsew signal input
flabel metal2 s 508784 -800 508896 480 0 FreeSans 1120 90 0 0 la_data_in[108]
port 173 nsew signal input
flabel metal2 s 512330 -800 512442 480 0 FreeSans 1120 90 0 0 la_data_in[109]
port 174 nsew signal input
flabel metal2 s 161276 -800 161388 480 0 FreeSans 1120 90 0 0 la_data_in[10]
port 175 nsew signal input
flabel metal2 s 515876 -800 515988 480 0 FreeSans 1120 90 0 0 la_data_in[110]
port 176 nsew signal input
flabel metal2 s 519422 -800 519534 480 0 FreeSans 1120 90 0 0 la_data_in[111]
port 177 nsew signal input
flabel metal2 s 522968 -800 523080 480 0 FreeSans 1120 90 0 0 la_data_in[112]
port 178 nsew signal input
flabel metal2 s 526514 -800 526626 480 0 FreeSans 1120 90 0 0 la_data_in[113]
port 179 nsew signal input
flabel metal2 s 530060 -800 530172 480 0 FreeSans 1120 90 0 0 la_data_in[114]
port 180 nsew signal input
flabel metal2 s 533606 -800 533718 480 0 FreeSans 1120 90 0 0 la_data_in[115]
port 181 nsew signal input
flabel metal2 s 537152 -800 537264 480 0 FreeSans 1120 90 0 0 la_data_in[116]
port 182 nsew signal input
flabel metal2 s 540698 -800 540810 480 0 FreeSans 1120 90 0 0 la_data_in[117]
port 183 nsew signal input
flabel metal2 s 544244 -800 544356 480 0 FreeSans 1120 90 0 0 la_data_in[118]
port 184 nsew signal input
flabel metal2 s 547790 -800 547902 480 0 FreeSans 1120 90 0 0 la_data_in[119]
port 185 nsew signal input
flabel metal2 s 164822 -800 164934 480 0 FreeSans 1120 90 0 0 la_data_in[11]
port 186 nsew signal input
flabel metal2 s 551336 -800 551448 480 0 FreeSans 1120 90 0 0 la_data_in[120]
port 187 nsew signal input
flabel metal2 s 554882 -800 554994 480 0 FreeSans 1120 90 0 0 la_data_in[121]
port 188 nsew signal input
flabel metal2 s 558428 -800 558540 480 0 FreeSans 1120 90 0 0 la_data_in[122]
port 189 nsew signal input
flabel metal2 s 561974 -800 562086 480 0 FreeSans 1120 90 0 0 la_data_in[123]
port 190 nsew signal input
flabel metal2 s 565520 -800 565632 480 0 FreeSans 1120 90 0 0 la_data_in[124]
port 191 nsew signal input
flabel metal2 s 569066 -800 569178 480 0 FreeSans 1120 90 0 0 la_data_in[125]
port 192 nsew signal input
flabel metal2 s 572612 -800 572724 480 0 FreeSans 1120 90 0 0 la_data_in[126]
port 193 nsew signal input
flabel metal2 s 576158 -800 576270 480 0 FreeSans 1120 90 0 0 la_data_in[127]
port 194 nsew signal input
flabel metal2 s 168368 -800 168480 480 0 FreeSans 1120 90 0 0 la_data_in[12]
port 195 nsew signal input
flabel metal2 s 171914 -800 172026 480 0 FreeSans 1120 90 0 0 la_data_in[13]
port 196 nsew signal input
flabel metal2 s 175460 -800 175572 480 0 FreeSans 1120 90 0 0 la_data_in[14]
port 197 nsew signal input
flabel metal2 s 179006 -800 179118 480 0 FreeSans 1120 90 0 0 la_data_in[15]
port 198 nsew signal input
flabel metal2 s 182552 -800 182664 480 0 FreeSans 1120 90 0 0 la_data_in[16]
port 199 nsew signal input
flabel metal2 s 186098 -800 186210 480 0 FreeSans 1120 90 0 0 la_data_in[17]
port 200 nsew signal input
flabel metal2 s 189644 -800 189756 480 0 FreeSans 1120 90 0 0 la_data_in[18]
port 201 nsew signal input
flabel metal2 s 193190 -800 193302 480 0 FreeSans 1120 90 0 0 la_data_in[19]
port 202 nsew signal input
flabel metal2 s 129362 -800 129474 480 0 FreeSans 1120 90 0 0 la_data_in[1]
port 203 nsew signal input
flabel metal2 s 196736 -800 196848 480 0 FreeSans 1120 90 0 0 la_data_in[20]
port 204 nsew signal input
flabel metal2 s 200282 -800 200394 480 0 FreeSans 1120 90 0 0 la_data_in[21]
port 205 nsew signal input
flabel metal2 s 203828 -800 203940 480 0 FreeSans 1120 90 0 0 la_data_in[22]
port 206 nsew signal input
flabel metal2 s 207374 -800 207486 480 0 FreeSans 1120 90 0 0 la_data_in[23]
port 207 nsew signal input
flabel metal2 s 210920 -800 211032 480 0 FreeSans 1120 90 0 0 la_data_in[24]
port 208 nsew signal input
flabel metal2 s 214466 -800 214578 480 0 FreeSans 1120 90 0 0 la_data_in[25]
port 209 nsew signal input
flabel metal2 s 218012 -800 218124 480 0 FreeSans 1120 90 0 0 la_data_in[26]
port 210 nsew signal input
flabel metal2 s 221558 -800 221670 480 0 FreeSans 1120 90 0 0 la_data_in[27]
port 211 nsew signal input
flabel metal2 s 225104 -800 225216 480 0 FreeSans 1120 90 0 0 la_data_in[28]
port 212 nsew signal input
flabel metal2 s 228650 -800 228762 480 0 FreeSans 1120 90 0 0 la_data_in[29]
port 213 nsew signal input
flabel metal2 s 132908 -800 133020 480 0 FreeSans 1120 90 0 0 la_data_in[2]
port 214 nsew signal input
flabel metal2 s 232196 -800 232308 480 0 FreeSans 1120 90 0 0 la_data_in[30]
port 215 nsew signal input
flabel metal2 s 235742 -800 235854 480 0 FreeSans 1120 90 0 0 la_data_in[31]
port 216 nsew signal input
flabel metal2 s 239288 -800 239400 480 0 FreeSans 1120 90 0 0 la_data_in[32]
port 217 nsew signal input
flabel metal2 s 242834 -800 242946 480 0 FreeSans 1120 90 0 0 la_data_in[33]
port 218 nsew signal input
flabel metal2 s 246380 -800 246492 480 0 FreeSans 1120 90 0 0 la_data_in[34]
port 219 nsew signal input
flabel metal2 s 249926 -800 250038 480 0 FreeSans 1120 90 0 0 la_data_in[35]
port 220 nsew signal input
flabel metal2 s 253472 -800 253584 480 0 FreeSans 1120 90 0 0 la_data_in[36]
port 221 nsew signal input
flabel metal2 s 257018 -800 257130 480 0 FreeSans 1120 90 0 0 la_data_in[37]
port 222 nsew signal input
flabel metal2 s 260564 -800 260676 480 0 FreeSans 1120 90 0 0 la_data_in[38]
port 223 nsew signal input
flabel metal2 s 264110 -800 264222 480 0 FreeSans 1120 90 0 0 la_data_in[39]
port 224 nsew signal input
flabel metal2 s 136454 -800 136566 480 0 FreeSans 1120 90 0 0 la_data_in[3]
port 225 nsew signal input
flabel metal2 s 267656 -800 267768 480 0 FreeSans 1120 90 0 0 la_data_in[40]
port 226 nsew signal input
flabel metal2 s 271202 -800 271314 480 0 FreeSans 1120 90 0 0 la_data_in[41]
port 227 nsew signal input
flabel metal2 s 274748 -800 274860 480 0 FreeSans 1120 90 0 0 la_data_in[42]
port 228 nsew signal input
flabel metal2 s 278294 -800 278406 480 0 FreeSans 1120 90 0 0 la_data_in[43]
port 229 nsew signal input
flabel metal2 s 281840 -800 281952 480 0 FreeSans 1120 90 0 0 la_data_in[44]
port 230 nsew signal input
flabel metal2 s 285386 -800 285498 480 0 FreeSans 1120 90 0 0 la_data_in[45]
port 231 nsew signal input
flabel metal2 s 288932 -800 289044 480 0 FreeSans 1120 90 0 0 la_data_in[46]
port 232 nsew signal input
flabel metal2 s 292478 -800 292590 480 0 FreeSans 1120 90 0 0 la_data_in[47]
port 233 nsew signal input
flabel metal2 s 296024 -800 296136 480 0 FreeSans 1120 90 0 0 la_data_in[48]
port 234 nsew signal input
flabel metal2 s 299570 -800 299682 480 0 FreeSans 1120 90 0 0 la_data_in[49]
port 235 nsew signal input
flabel metal2 s 140000 -800 140112 480 0 FreeSans 1120 90 0 0 la_data_in[4]
port 236 nsew signal input
flabel metal2 s 303116 -800 303228 480 0 FreeSans 1120 90 0 0 la_data_in[50]
port 237 nsew signal input
flabel metal2 s 306662 -800 306774 480 0 FreeSans 1120 90 0 0 la_data_in[51]
port 238 nsew signal input
flabel metal2 s 310208 -800 310320 480 0 FreeSans 1120 90 0 0 la_data_in[52]
port 239 nsew signal input
flabel metal2 s 313754 -800 313866 480 0 FreeSans 1120 90 0 0 la_data_in[53]
port 240 nsew signal input
flabel metal2 s 317300 -800 317412 480 0 FreeSans 1120 90 0 0 la_data_in[54]
port 241 nsew signal input
flabel metal2 s 320846 -800 320958 480 0 FreeSans 1120 90 0 0 la_data_in[55]
port 242 nsew signal input
flabel metal2 s 324392 -800 324504 480 0 FreeSans 1120 90 0 0 la_data_in[56]
port 243 nsew signal input
flabel metal2 s 327938 -800 328050 480 0 FreeSans 1120 90 0 0 la_data_in[57]
port 244 nsew signal input
flabel metal2 s 331484 -800 331596 480 0 FreeSans 1120 90 0 0 la_data_in[58]
port 245 nsew signal input
flabel metal2 s 335030 -800 335142 480 0 FreeSans 1120 90 0 0 la_data_in[59]
port 246 nsew signal input
flabel metal2 s 143546 -800 143658 480 0 FreeSans 1120 90 0 0 la_data_in[5]
port 247 nsew signal input
flabel metal2 s 338576 -800 338688 480 0 FreeSans 1120 90 0 0 la_data_in[60]
port 248 nsew signal input
flabel metal2 s 342122 -800 342234 480 0 FreeSans 1120 90 0 0 la_data_in[61]
port 249 nsew signal input
flabel metal2 s 345668 -800 345780 480 0 FreeSans 1120 90 0 0 la_data_in[62]
port 250 nsew signal input
flabel metal2 s 349214 -800 349326 480 0 FreeSans 1120 90 0 0 la_data_in[63]
port 251 nsew signal input
flabel metal2 s 352760 -800 352872 480 0 FreeSans 1120 90 0 0 la_data_in[64]
port 252 nsew signal input
flabel metal2 s 356306 -800 356418 480 0 FreeSans 1120 90 0 0 la_data_in[65]
port 253 nsew signal input
flabel metal2 s 359852 -800 359964 480 0 FreeSans 1120 90 0 0 la_data_in[66]
port 254 nsew signal input
flabel metal2 s 363398 -800 363510 480 0 FreeSans 1120 90 0 0 la_data_in[67]
port 255 nsew signal input
flabel metal2 s 366944 -800 367056 480 0 FreeSans 1120 90 0 0 la_data_in[68]
port 256 nsew signal input
flabel metal2 s 370490 -800 370602 480 0 FreeSans 1120 90 0 0 la_data_in[69]
port 257 nsew signal input
flabel metal2 s 147092 -800 147204 480 0 FreeSans 1120 90 0 0 la_data_in[6]
port 258 nsew signal input
flabel metal2 s 374036 -800 374148 480 0 FreeSans 1120 90 0 0 la_data_in[70]
port 259 nsew signal input
flabel metal2 s 377582 -800 377694 480 0 FreeSans 1120 90 0 0 la_data_in[71]
port 260 nsew signal input
flabel metal2 s 381128 -800 381240 480 0 FreeSans 1120 90 0 0 la_data_in[72]
port 261 nsew signal input
flabel metal2 s 384674 -800 384786 480 0 FreeSans 1120 90 0 0 la_data_in[73]
port 262 nsew signal input
flabel metal2 s 388220 -800 388332 480 0 FreeSans 1120 90 0 0 la_data_in[74]
port 263 nsew signal input
flabel metal2 s 391766 -800 391878 480 0 FreeSans 1120 90 0 0 la_data_in[75]
port 264 nsew signal input
flabel metal2 s 395312 -800 395424 480 0 FreeSans 1120 90 0 0 la_data_in[76]
port 265 nsew signal input
flabel metal2 s 398858 -800 398970 480 0 FreeSans 1120 90 0 0 la_data_in[77]
port 266 nsew signal input
flabel metal2 s 402404 -800 402516 480 0 FreeSans 1120 90 0 0 la_data_in[78]
port 267 nsew signal input
flabel metal2 s 405950 -800 406062 480 0 FreeSans 1120 90 0 0 la_data_in[79]
port 268 nsew signal input
flabel metal2 s 150638 -800 150750 480 0 FreeSans 1120 90 0 0 la_data_in[7]
port 269 nsew signal input
flabel metal2 s 409496 -800 409608 480 0 FreeSans 1120 90 0 0 la_data_in[80]
port 270 nsew signal input
flabel metal2 s 413042 -800 413154 480 0 FreeSans 1120 90 0 0 la_data_in[81]
port 271 nsew signal input
flabel metal2 s 416588 -800 416700 480 0 FreeSans 1120 90 0 0 la_data_in[82]
port 272 nsew signal input
flabel metal2 s 420134 -800 420246 480 0 FreeSans 1120 90 0 0 la_data_in[83]
port 273 nsew signal input
flabel metal2 s 423680 -800 423792 480 0 FreeSans 1120 90 0 0 la_data_in[84]
port 274 nsew signal input
flabel metal2 s 427226 -800 427338 480 0 FreeSans 1120 90 0 0 la_data_in[85]
port 275 nsew signal input
flabel metal2 s 430772 -800 430884 480 0 FreeSans 1120 90 0 0 la_data_in[86]
port 276 nsew signal input
flabel metal2 s 434318 -800 434430 480 0 FreeSans 1120 90 0 0 la_data_in[87]
port 277 nsew signal input
flabel metal2 s 437864 -800 437976 480 0 FreeSans 1120 90 0 0 la_data_in[88]
port 278 nsew signal input
flabel metal2 s 441410 -800 441522 480 0 FreeSans 1120 90 0 0 la_data_in[89]
port 279 nsew signal input
flabel metal2 s 154184 -800 154296 480 0 FreeSans 1120 90 0 0 la_data_in[8]
port 280 nsew signal input
flabel metal2 s 444956 -800 445068 480 0 FreeSans 1120 90 0 0 la_data_in[90]
port 281 nsew signal input
flabel metal2 s 448502 -800 448614 480 0 FreeSans 1120 90 0 0 la_data_in[91]
port 282 nsew signal input
flabel metal2 s 452048 -800 452160 480 0 FreeSans 1120 90 0 0 la_data_in[92]
port 283 nsew signal input
flabel metal2 s 455594 -800 455706 480 0 FreeSans 1120 90 0 0 la_data_in[93]
port 284 nsew signal input
flabel metal2 s 459140 -800 459252 480 0 FreeSans 1120 90 0 0 la_data_in[94]
port 285 nsew signal input
flabel metal2 s 462686 -800 462798 480 0 FreeSans 1120 90 0 0 la_data_in[95]
port 286 nsew signal input
flabel metal2 s 466232 -800 466344 480 0 FreeSans 1120 90 0 0 la_data_in[96]
port 287 nsew signal input
flabel metal2 s 469778 -800 469890 480 0 FreeSans 1120 90 0 0 la_data_in[97]
port 288 nsew signal input
flabel metal2 s 473324 -800 473436 480 0 FreeSans 1120 90 0 0 la_data_in[98]
port 289 nsew signal input
flabel metal2 s 476870 -800 476982 480 0 FreeSans 1120 90 0 0 la_data_in[99]
port 290 nsew signal input
flabel metal2 s 157730 -800 157842 480 0 FreeSans 1120 90 0 0 la_data_in[9]
port 291 nsew signal input
flabel metal2 s 126998 -800 127110 480 0 FreeSans 1120 90 0 0 la_data_out[0]
port 292 nsew signal tristate
flabel metal2 s 481598 -800 481710 480 0 FreeSans 1120 90 0 0 la_data_out[100]
port 293 nsew signal tristate
flabel metal2 s 485144 -800 485256 480 0 FreeSans 1120 90 0 0 la_data_out[101]
port 294 nsew signal tristate
flabel metal2 s 488690 -800 488802 480 0 FreeSans 1120 90 0 0 la_data_out[102]
port 295 nsew signal tristate
flabel metal2 s 492236 -800 492348 480 0 FreeSans 1120 90 0 0 la_data_out[103]
port 296 nsew signal tristate
flabel metal2 s 495782 -800 495894 480 0 FreeSans 1120 90 0 0 la_data_out[104]
port 297 nsew signal tristate
flabel metal2 s 499328 -800 499440 480 0 FreeSans 1120 90 0 0 la_data_out[105]
port 298 nsew signal tristate
flabel metal2 s 502874 -800 502986 480 0 FreeSans 1120 90 0 0 la_data_out[106]
port 299 nsew signal tristate
flabel metal2 s 506420 -800 506532 480 0 FreeSans 1120 90 0 0 la_data_out[107]
port 300 nsew signal tristate
flabel metal2 s 509966 -800 510078 480 0 FreeSans 1120 90 0 0 la_data_out[108]
port 301 nsew signal tristate
flabel metal2 s 513512 -800 513624 480 0 FreeSans 1120 90 0 0 la_data_out[109]
port 302 nsew signal tristate
flabel metal2 s 162458 -800 162570 480 0 FreeSans 1120 90 0 0 la_data_out[10]
port 303 nsew signal tristate
flabel metal2 s 517058 -800 517170 480 0 FreeSans 1120 90 0 0 la_data_out[110]
port 304 nsew signal tristate
flabel metal2 s 520604 -800 520716 480 0 FreeSans 1120 90 0 0 la_data_out[111]
port 305 nsew signal tristate
flabel metal2 s 524150 -800 524262 480 0 FreeSans 1120 90 0 0 la_data_out[112]
port 306 nsew signal tristate
flabel metal2 s 527696 -800 527808 480 0 FreeSans 1120 90 0 0 la_data_out[113]
port 307 nsew signal tristate
flabel metal2 s 531242 -800 531354 480 0 FreeSans 1120 90 0 0 la_data_out[114]
port 308 nsew signal tristate
flabel metal2 s 534788 -800 534900 480 0 FreeSans 1120 90 0 0 la_data_out[115]
port 309 nsew signal tristate
flabel metal2 s 538334 -800 538446 480 0 FreeSans 1120 90 0 0 la_data_out[116]
port 310 nsew signal tristate
flabel metal2 s 541880 -800 541992 480 0 FreeSans 1120 90 0 0 la_data_out[117]
port 311 nsew signal tristate
flabel metal2 s 545426 -800 545538 480 0 FreeSans 1120 90 0 0 la_data_out[118]
port 312 nsew signal tristate
flabel metal2 s 548972 -800 549084 480 0 FreeSans 1120 90 0 0 la_data_out[119]
port 313 nsew signal tristate
flabel metal2 s 166004 -800 166116 480 0 FreeSans 1120 90 0 0 la_data_out[11]
port 314 nsew signal tristate
flabel metal2 s 552518 -800 552630 480 0 FreeSans 1120 90 0 0 la_data_out[120]
port 315 nsew signal tristate
flabel metal2 s 556064 -800 556176 480 0 FreeSans 1120 90 0 0 la_data_out[121]
port 316 nsew signal tristate
flabel metal2 s 559610 -800 559722 480 0 FreeSans 1120 90 0 0 la_data_out[122]
port 317 nsew signal tristate
flabel metal2 s 563156 -800 563268 480 0 FreeSans 1120 90 0 0 la_data_out[123]
port 318 nsew signal tristate
flabel metal2 s 566702 -800 566814 480 0 FreeSans 1120 90 0 0 la_data_out[124]
port 319 nsew signal tristate
flabel metal2 s 570248 -800 570360 480 0 FreeSans 1120 90 0 0 la_data_out[125]
port 320 nsew signal tristate
flabel metal2 s 573794 -800 573906 480 0 FreeSans 1120 90 0 0 la_data_out[126]
port 321 nsew signal tristate
flabel metal2 s 577340 -800 577452 480 0 FreeSans 1120 90 0 0 la_data_out[127]
port 322 nsew signal tristate
flabel metal2 s 169550 -800 169662 480 0 FreeSans 1120 90 0 0 la_data_out[12]
port 323 nsew signal tristate
flabel metal2 s 173096 -800 173208 480 0 FreeSans 1120 90 0 0 la_data_out[13]
port 324 nsew signal tristate
flabel metal2 s 176642 -800 176754 480 0 FreeSans 1120 90 0 0 la_data_out[14]
port 325 nsew signal tristate
flabel metal2 s 180188 -800 180300 480 0 FreeSans 1120 90 0 0 la_data_out[15]
port 326 nsew signal tristate
flabel metal2 s 183734 -800 183846 480 0 FreeSans 1120 90 0 0 la_data_out[16]
port 327 nsew signal tristate
flabel metal2 s 187280 -800 187392 480 0 FreeSans 1120 90 0 0 la_data_out[17]
port 328 nsew signal tristate
flabel metal2 s 190826 -800 190938 480 0 FreeSans 1120 90 0 0 la_data_out[18]
port 329 nsew signal tristate
flabel metal2 s 194372 -800 194484 480 0 FreeSans 1120 90 0 0 la_data_out[19]
port 330 nsew signal tristate
flabel metal2 s 130544 -800 130656 480 0 FreeSans 1120 90 0 0 la_data_out[1]
port 331 nsew signal tristate
flabel metal2 s 197918 -800 198030 480 0 FreeSans 1120 90 0 0 la_data_out[20]
port 332 nsew signal tristate
flabel metal2 s 201464 -800 201576 480 0 FreeSans 1120 90 0 0 la_data_out[21]
port 333 nsew signal tristate
flabel metal2 s 205010 -800 205122 480 0 FreeSans 1120 90 0 0 la_data_out[22]
port 334 nsew signal tristate
flabel metal2 s 208556 -800 208668 480 0 FreeSans 1120 90 0 0 la_data_out[23]
port 335 nsew signal tristate
flabel metal2 s 212102 -800 212214 480 0 FreeSans 1120 90 0 0 la_data_out[24]
port 336 nsew signal tristate
flabel metal2 s 215648 -800 215760 480 0 FreeSans 1120 90 0 0 la_data_out[25]
port 337 nsew signal tristate
flabel metal2 s 219194 -800 219306 480 0 FreeSans 1120 90 0 0 la_data_out[26]
port 338 nsew signal tristate
flabel metal2 s 222740 -800 222852 480 0 FreeSans 1120 90 0 0 la_data_out[27]
port 339 nsew signal tristate
flabel metal2 s 226286 -800 226398 480 0 FreeSans 1120 90 0 0 la_data_out[28]
port 340 nsew signal tristate
flabel metal2 s 229832 -800 229944 480 0 FreeSans 1120 90 0 0 la_data_out[29]
port 341 nsew signal tristate
flabel metal2 s 134090 -800 134202 480 0 FreeSans 1120 90 0 0 la_data_out[2]
port 342 nsew signal tristate
flabel metal2 s 233378 -800 233490 480 0 FreeSans 1120 90 0 0 la_data_out[30]
port 343 nsew signal tristate
flabel metal2 s 236924 -800 237036 480 0 FreeSans 1120 90 0 0 la_data_out[31]
port 344 nsew signal tristate
flabel metal2 s 240470 -800 240582 480 0 FreeSans 1120 90 0 0 la_data_out[32]
port 345 nsew signal tristate
flabel metal2 s 244016 -800 244128 480 0 FreeSans 1120 90 0 0 la_data_out[33]
port 346 nsew signal tristate
flabel metal2 s 247562 -800 247674 480 0 FreeSans 1120 90 0 0 la_data_out[34]
port 347 nsew signal tristate
flabel metal2 s 251108 -800 251220 480 0 FreeSans 1120 90 0 0 la_data_out[35]
port 348 nsew signal tristate
flabel metal2 s 254654 -800 254766 480 0 FreeSans 1120 90 0 0 la_data_out[36]
port 349 nsew signal tristate
flabel metal2 s 258200 -800 258312 480 0 FreeSans 1120 90 0 0 la_data_out[37]
port 350 nsew signal tristate
flabel metal2 s 261746 -800 261858 480 0 FreeSans 1120 90 0 0 la_data_out[38]
port 351 nsew signal tristate
flabel metal2 s 265292 -800 265404 480 0 FreeSans 1120 90 0 0 la_data_out[39]
port 352 nsew signal tristate
flabel metal2 s 137636 -800 137748 480 0 FreeSans 1120 90 0 0 la_data_out[3]
port 353 nsew signal tristate
flabel metal2 s 268838 -800 268950 480 0 FreeSans 1120 90 0 0 la_data_out[40]
port 354 nsew signal tristate
flabel metal2 s 272384 -800 272496 480 0 FreeSans 1120 90 0 0 la_data_out[41]
port 355 nsew signal tristate
flabel metal2 s 275930 -800 276042 480 0 FreeSans 1120 90 0 0 la_data_out[42]
port 356 nsew signal tristate
flabel metal2 s 279476 -800 279588 480 0 FreeSans 1120 90 0 0 la_data_out[43]
port 357 nsew signal tristate
flabel metal2 s 283022 -800 283134 480 0 FreeSans 1120 90 0 0 la_data_out[44]
port 358 nsew signal tristate
flabel metal2 s 286568 -800 286680 480 0 FreeSans 1120 90 0 0 la_data_out[45]
port 359 nsew signal tristate
flabel metal2 s 290114 -800 290226 480 0 FreeSans 1120 90 0 0 la_data_out[46]
port 360 nsew signal tristate
flabel metal2 s 293660 -800 293772 480 0 FreeSans 1120 90 0 0 la_data_out[47]
port 361 nsew signal tristate
flabel metal2 s 297206 -800 297318 480 0 FreeSans 1120 90 0 0 la_data_out[48]
port 362 nsew signal tristate
flabel metal2 s 300752 -800 300864 480 0 FreeSans 1120 90 0 0 la_data_out[49]
port 363 nsew signal tristate
flabel metal2 s 141182 -800 141294 480 0 FreeSans 1120 90 0 0 la_data_out[4]
port 364 nsew signal tristate
flabel metal2 s 304298 -800 304410 480 0 FreeSans 1120 90 0 0 la_data_out[50]
port 365 nsew signal tristate
flabel metal2 s 307844 -800 307956 480 0 FreeSans 1120 90 0 0 la_data_out[51]
port 366 nsew signal tristate
flabel metal2 s 311390 -800 311502 480 0 FreeSans 1120 90 0 0 la_data_out[52]
port 367 nsew signal tristate
flabel metal2 s 314936 -800 315048 480 0 FreeSans 1120 90 0 0 la_data_out[53]
port 368 nsew signal tristate
flabel metal2 s 318482 -800 318594 480 0 FreeSans 1120 90 0 0 la_data_out[54]
port 369 nsew signal tristate
flabel metal2 s 322028 -800 322140 480 0 FreeSans 1120 90 0 0 la_data_out[55]
port 370 nsew signal tristate
flabel metal2 s 325574 -800 325686 480 0 FreeSans 1120 90 0 0 la_data_out[56]
port 371 nsew signal tristate
flabel metal2 s 329120 -800 329232 480 0 FreeSans 1120 90 0 0 la_data_out[57]
port 372 nsew signal tristate
flabel metal2 s 332666 -800 332778 480 0 FreeSans 1120 90 0 0 la_data_out[58]
port 373 nsew signal tristate
flabel metal2 s 336212 -800 336324 480 0 FreeSans 1120 90 0 0 la_data_out[59]
port 374 nsew signal tristate
flabel metal2 s 144728 -800 144840 480 0 FreeSans 1120 90 0 0 la_data_out[5]
port 375 nsew signal tristate
flabel metal2 s 339758 -800 339870 480 0 FreeSans 1120 90 0 0 la_data_out[60]
port 376 nsew signal tristate
flabel metal2 s 343304 -800 343416 480 0 FreeSans 1120 90 0 0 la_data_out[61]
port 377 nsew signal tristate
flabel metal2 s 346850 -800 346962 480 0 FreeSans 1120 90 0 0 la_data_out[62]
port 378 nsew signal tristate
flabel metal2 s 350396 -800 350508 480 0 FreeSans 1120 90 0 0 la_data_out[63]
port 379 nsew signal tristate
flabel metal2 s 353942 -800 354054 480 0 FreeSans 1120 90 0 0 la_data_out[64]
port 380 nsew signal tristate
flabel metal2 s 357488 -800 357600 480 0 FreeSans 1120 90 0 0 la_data_out[65]
port 381 nsew signal tristate
flabel metal2 s 361034 -800 361146 480 0 FreeSans 1120 90 0 0 la_data_out[66]
port 382 nsew signal tristate
flabel metal2 s 364580 -800 364692 480 0 FreeSans 1120 90 0 0 la_data_out[67]
port 383 nsew signal tristate
flabel metal2 s 368126 -800 368238 480 0 FreeSans 1120 90 0 0 la_data_out[68]
port 384 nsew signal tristate
flabel metal2 s 371672 -800 371784 480 0 FreeSans 1120 90 0 0 la_data_out[69]
port 385 nsew signal tristate
flabel metal2 s 148274 -800 148386 480 0 FreeSans 1120 90 0 0 la_data_out[6]
port 386 nsew signal tristate
flabel metal2 s 375218 -800 375330 480 0 FreeSans 1120 90 0 0 la_data_out[70]
port 387 nsew signal tristate
flabel metal2 s 378764 -800 378876 480 0 FreeSans 1120 90 0 0 la_data_out[71]
port 388 nsew signal tristate
flabel metal2 s 382310 -800 382422 480 0 FreeSans 1120 90 0 0 la_data_out[72]
port 389 nsew signal tristate
flabel metal2 s 385856 -800 385968 480 0 FreeSans 1120 90 0 0 la_data_out[73]
port 390 nsew signal tristate
flabel metal2 s 389402 -800 389514 480 0 FreeSans 1120 90 0 0 la_data_out[74]
port 391 nsew signal tristate
flabel metal2 s 392948 -800 393060 480 0 FreeSans 1120 90 0 0 la_data_out[75]
port 392 nsew signal tristate
flabel metal2 s 396494 -800 396606 480 0 FreeSans 1120 90 0 0 la_data_out[76]
port 393 nsew signal tristate
flabel metal2 s 400040 -800 400152 480 0 FreeSans 1120 90 0 0 la_data_out[77]
port 394 nsew signal tristate
flabel metal2 s 403586 -800 403698 480 0 FreeSans 1120 90 0 0 la_data_out[78]
port 395 nsew signal tristate
flabel metal2 s 407132 -800 407244 480 0 FreeSans 1120 90 0 0 la_data_out[79]
port 396 nsew signal tristate
flabel metal2 s 151820 -800 151932 480 0 FreeSans 1120 90 0 0 la_data_out[7]
port 397 nsew signal tristate
flabel metal2 s 410678 -800 410790 480 0 FreeSans 1120 90 0 0 la_data_out[80]
port 398 nsew signal tristate
flabel metal2 s 414224 -800 414336 480 0 FreeSans 1120 90 0 0 la_data_out[81]
port 399 nsew signal tristate
flabel metal2 s 417770 -800 417882 480 0 FreeSans 1120 90 0 0 la_data_out[82]
port 400 nsew signal tristate
flabel metal2 s 421316 -800 421428 480 0 FreeSans 1120 90 0 0 la_data_out[83]
port 401 nsew signal tristate
flabel metal2 s 424862 -800 424974 480 0 FreeSans 1120 90 0 0 la_data_out[84]
port 402 nsew signal tristate
flabel metal2 s 428408 -800 428520 480 0 FreeSans 1120 90 0 0 la_data_out[85]
port 403 nsew signal tristate
flabel metal2 s 431954 -800 432066 480 0 FreeSans 1120 90 0 0 la_data_out[86]
port 404 nsew signal tristate
flabel metal2 s 435500 -800 435612 480 0 FreeSans 1120 90 0 0 la_data_out[87]
port 405 nsew signal tristate
flabel metal2 s 439046 -800 439158 480 0 FreeSans 1120 90 0 0 la_data_out[88]
port 406 nsew signal tristate
flabel metal2 s 442592 -800 442704 480 0 FreeSans 1120 90 0 0 la_data_out[89]
port 407 nsew signal tristate
flabel metal2 s 155366 -800 155478 480 0 FreeSans 1120 90 0 0 la_data_out[8]
port 408 nsew signal tristate
flabel metal2 s 446138 -800 446250 480 0 FreeSans 1120 90 0 0 la_data_out[90]
port 409 nsew signal tristate
flabel metal2 s 449684 -800 449796 480 0 FreeSans 1120 90 0 0 la_data_out[91]
port 410 nsew signal tristate
flabel metal2 s 453230 -800 453342 480 0 FreeSans 1120 90 0 0 la_data_out[92]
port 411 nsew signal tristate
flabel metal2 s 456776 -800 456888 480 0 FreeSans 1120 90 0 0 la_data_out[93]
port 412 nsew signal tristate
flabel metal2 s 460322 -800 460434 480 0 FreeSans 1120 90 0 0 la_data_out[94]
port 413 nsew signal tristate
flabel metal2 s 463868 -800 463980 480 0 FreeSans 1120 90 0 0 la_data_out[95]
port 414 nsew signal tristate
flabel metal2 s 467414 -800 467526 480 0 FreeSans 1120 90 0 0 la_data_out[96]
port 415 nsew signal tristate
flabel metal2 s 470960 -800 471072 480 0 FreeSans 1120 90 0 0 la_data_out[97]
port 416 nsew signal tristate
flabel metal2 s 474506 -800 474618 480 0 FreeSans 1120 90 0 0 la_data_out[98]
port 417 nsew signal tristate
flabel metal2 s 478052 -800 478164 480 0 FreeSans 1120 90 0 0 la_data_out[99]
port 418 nsew signal tristate
flabel metal2 s 158912 -800 159024 480 0 FreeSans 1120 90 0 0 la_data_out[9]
port 419 nsew signal tristate
flabel metal2 s 128180 -800 128292 480 0 FreeSans 1120 90 0 0 la_oenb[0]
port 420 nsew signal input
flabel metal2 s 482780 -800 482892 480 0 FreeSans 1120 90 0 0 la_oenb[100]
port 421 nsew signal input
flabel metal2 s 486326 -800 486438 480 0 FreeSans 1120 90 0 0 la_oenb[101]
port 422 nsew signal input
flabel metal2 s 489872 -800 489984 480 0 FreeSans 1120 90 0 0 la_oenb[102]
port 423 nsew signal input
flabel metal2 s 493418 -800 493530 480 0 FreeSans 1120 90 0 0 la_oenb[103]
port 424 nsew signal input
flabel metal2 s 496964 -800 497076 480 0 FreeSans 1120 90 0 0 la_oenb[104]
port 425 nsew signal input
flabel metal2 s 500510 -800 500622 480 0 FreeSans 1120 90 0 0 la_oenb[105]
port 426 nsew signal input
flabel metal2 s 504056 -800 504168 480 0 FreeSans 1120 90 0 0 la_oenb[106]
port 427 nsew signal input
flabel metal2 s 507602 -800 507714 480 0 FreeSans 1120 90 0 0 la_oenb[107]
port 428 nsew signal input
flabel metal2 s 511148 -800 511260 480 0 FreeSans 1120 90 0 0 la_oenb[108]
port 429 nsew signal input
flabel metal2 s 514694 -800 514806 480 0 FreeSans 1120 90 0 0 la_oenb[109]
port 430 nsew signal input
flabel metal2 s 163640 -800 163752 480 0 FreeSans 1120 90 0 0 la_oenb[10]
port 431 nsew signal input
flabel metal2 s 518240 -800 518352 480 0 FreeSans 1120 90 0 0 la_oenb[110]
port 432 nsew signal input
flabel metal2 s 521786 -800 521898 480 0 FreeSans 1120 90 0 0 la_oenb[111]
port 433 nsew signal input
flabel metal2 s 525332 -800 525444 480 0 FreeSans 1120 90 0 0 la_oenb[112]
port 434 nsew signal input
flabel metal2 s 528878 -800 528990 480 0 FreeSans 1120 90 0 0 la_oenb[113]
port 435 nsew signal input
flabel metal2 s 532424 -800 532536 480 0 FreeSans 1120 90 0 0 la_oenb[114]
port 436 nsew signal input
flabel metal2 s 535970 -800 536082 480 0 FreeSans 1120 90 0 0 la_oenb[115]
port 437 nsew signal input
flabel metal2 s 539516 -800 539628 480 0 FreeSans 1120 90 0 0 la_oenb[116]
port 438 nsew signal input
flabel metal2 s 543062 -800 543174 480 0 FreeSans 1120 90 0 0 la_oenb[117]
port 439 nsew signal input
flabel metal2 s 546608 -800 546720 480 0 FreeSans 1120 90 0 0 la_oenb[118]
port 440 nsew signal input
flabel metal2 s 550154 -800 550266 480 0 FreeSans 1120 90 0 0 la_oenb[119]
port 441 nsew signal input
flabel metal2 s 167186 -800 167298 480 0 FreeSans 1120 90 0 0 la_oenb[11]
port 442 nsew signal input
flabel metal2 s 553700 -800 553812 480 0 FreeSans 1120 90 0 0 la_oenb[120]
port 443 nsew signal input
flabel metal2 s 557246 -800 557358 480 0 FreeSans 1120 90 0 0 la_oenb[121]
port 444 nsew signal input
flabel metal2 s 560792 -800 560904 480 0 FreeSans 1120 90 0 0 la_oenb[122]
port 445 nsew signal input
flabel metal2 s 564338 -800 564450 480 0 FreeSans 1120 90 0 0 la_oenb[123]
port 446 nsew signal input
flabel metal2 s 567884 -800 567996 480 0 FreeSans 1120 90 0 0 la_oenb[124]
port 447 nsew signal input
flabel metal2 s 571430 -800 571542 480 0 FreeSans 1120 90 0 0 la_oenb[125]
port 448 nsew signal input
flabel metal2 s 574976 -800 575088 480 0 FreeSans 1120 90 0 0 la_oenb[126]
port 449 nsew signal input
flabel metal2 s 578522 -800 578634 480 0 FreeSans 1120 90 0 0 la_oenb[127]
port 450 nsew signal input
flabel metal2 s 170732 -800 170844 480 0 FreeSans 1120 90 0 0 la_oenb[12]
port 451 nsew signal input
flabel metal2 s 174278 -800 174390 480 0 FreeSans 1120 90 0 0 la_oenb[13]
port 452 nsew signal input
flabel metal2 s 177824 -800 177936 480 0 FreeSans 1120 90 0 0 la_oenb[14]
port 453 nsew signal input
flabel metal2 s 181370 -800 181482 480 0 FreeSans 1120 90 0 0 la_oenb[15]
port 454 nsew signal input
flabel metal2 s 184916 -800 185028 480 0 FreeSans 1120 90 0 0 la_oenb[16]
port 455 nsew signal input
flabel metal2 s 188462 -800 188574 480 0 FreeSans 1120 90 0 0 la_oenb[17]
port 456 nsew signal input
flabel metal2 s 192008 -800 192120 480 0 FreeSans 1120 90 0 0 la_oenb[18]
port 457 nsew signal input
flabel metal2 s 195554 -800 195666 480 0 FreeSans 1120 90 0 0 la_oenb[19]
port 458 nsew signal input
flabel metal2 s 131726 -800 131838 480 0 FreeSans 1120 90 0 0 la_oenb[1]
port 459 nsew signal input
flabel metal2 s 199100 -800 199212 480 0 FreeSans 1120 90 0 0 la_oenb[20]
port 460 nsew signal input
flabel metal2 s 202646 -800 202758 480 0 FreeSans 1120 90 0 0 la_oenb[21]
port 461 nsew signal input
flabel metal2 s 206192 -800 206304 480 0 FreeSans 1120 90 0 0 la_oenb[22]
port 462 nsew signal input
flabel metal2 s 209738 -800 209850 480 0 FreeSans 1120 90 0 0 la_oenb[23]
port 463 nsew signal input
flabel metal2 s 213284 -800 213396 480 0 FreeSans 1120 90 0 0 la_oenb[24]
port 464 nsew signal input
flabel metal2 s 216830 -800 216942 480 0 FreeSans 1120 90 0 0 la_oenb[25]
port 465 nsew signal input
flabel metal2 s 220376 -800 220488 480 0 FreeSans 1120 90 0 0 la_oenb[26]
port 466 nsew signal input
flabel metal2 s 223922 -800 224034 480 0 FreeSans 1120 90 0 0 la_oenb[27]
port 467 nsew signal input
flabel metal2 s 227468 -800 227580 480 0 FreeSans 1120 90 0 0 la_oenb[28]
port 468 nsew signal input
flabel metal2 s 231014 -800 231126 480 0 FreeSans 1120 90 0 0 la_oenb[29]
port 469 nsew signal input
flabel metal2 s 135272 -800 135384 480 0 FreeSans 1120 90 0 0 la_oenb[2]
port 470 nsew signal input
flabel metal2 s 234560 -800 234672 480 0 FreeSans 1120 90 0 0 la_oenb[30]
port 471 nsew signal input
flabel metal2 s 238106 -800 238218 480 0 FreeSans 1120 90 0 0 la_oenb[31]
port 472 nsew signal input
flabel metal2 s 241652 -800 241764 480 0 FreeSans 1120 90 0 0 la_oenb[32]
port 473 nsew signal input
flabel metal2 s 245198 -800 245310 480 0 FreeSans 1120 90 0 0 la_oenb[33]
port 474 nsew signal input
flabel metal2 s 248744 -800 248856 480 0 FreeSans 1120 90 0 0 la_oenb[34]
port 475 nsew signal input
flabel metal2 s 252290 -800 252402 480 0 FreeSans 1120 90 0 0 la_oenb[35]
port 476 nsew signal input
flabel metal2 s 255836 -800 255948 480 0 FreeSans 1120 90 0 0 la_oenb[36]
port 477 nsew signal input
flabel metal2 s 259382 -800 259494 480 0 FreeSans 1120 90 0 0 la_oenb[37]
port 478 nsew signal input
flabel metal2 s 262928 -800 263040 480 0 FreeSans 1120 90 0 0 la_oenb[38]
port 479 nsew signal input
flabel metal2 s 266474 -800 266586 480 0 FreeSans 1120 90 0 0 la_oenb[39]
port 480 nsew signal input
flabel metal2 s 138818 -800 138930 480 0 FreeSans 1120 90 0 0 la_oenb[3]
port 481 nsew signal input
flabel metal2 s 270020 -800 270132 480 0 FreeSans 1120 90 0 0 la_oenb[40]
port 482 nsew signal input
flabel metal2 s 273566 -800 273678 480 0 FreeSans 1120 90 0 0 la_oenb[41]
port 483 nsew signal input
flabel metal2 s 277112 -800 277224 480 0 FreeSans 1120 90 0 0 la_oenb[42]
port 484 nsew signal input
flabel metal2 s 280658 -800 280770 480 0 FreeSans 1120 90 0 0 la_oenb[43]
port 485 nsew signal input
flabel metal2 s 284204 -800 284316 480 0 FreeSans 1120 90 0 0 la_oenb[44]
port 486 nsew signal input
flabel metal2 s 287750 -800 287862 480 0 FreeSans 1120 90 0 0 la_oenb[45]
port 487 nsew signal input
flabel metal2 s 291296 -800 291408 480 0 FreeSans 1120 90 0 0 la_oenb[46]
port 488 nsew signal input
flabel metal2 s 294842 -800 294954 480 0 FreeSans 1120 90 0 0 la_oenb[47]
port 489 nsew signal input
flabel metal2 s 298388 -800 298500 480 0 FreeSans 1120 90 0 0 la_oenb[48]
port 490 nsew signal input
flabel metal2 s 301934 -800 302046 480 0 FreeSans 1120 90 0 0 la_oenb[49]
port 491 nsew signal input
flabel metal2 s 142364 -800 142476 480 0 FreeSans 1120 90 0 0 la_oenb[4]
port 492 nsew signal input
flabel metal2 s 305480 -800 305592 480 0 FreeSans 1120 90 0 0 la_oenb[50]
port 493 nsew signal input
flabel metal2 s 309026 -800 309138 480 0 FreeSans 1120 90 0 0 la_oenb[51]
port 494 nsew signal input
flabel metal2 s 312572 -800 312684 480 0 FreeSans 1120 90 0 0 la_oenb[52]
port 495 nsew signal input
flabel metal2 s 316118 -800 316230 480 0 FreeSans 1120 90 0 0 la_oenb[53]
port 496 nsew signal input
flabel metal2 s 319664 -800 319776 480 0 FreeSans 1120 90 0 0 la_oenb[54]
port 497 nsew signal input
flabel metal2 s 323210 -800 323322 480 0 FreeSans 1120 90 0 0 la_oenb[55]
port 498 nsew signal input
flabel metal2 s 326756 -800 326868 480 0 FreeSans 1120 90 0 0 la_oenb[56]
port 499 nsew signal input
flabel metal2 s 330302 -800 330414 480 0 FreeSans 1120 90 0 0 la_oenb[57]
port 500 nsew signal input
flabel metal2 s 333848 -800 333960 480 0 FreeSans 1120 90 0 0 la_oenb[58]
port 501 nsew signal input
flabel metal2 s 337394 -800 337506 480 0 FreeSans 1120 90 0 0 la_oenb[59]
port 502 nsew signal input
flabel metal2 s 145910 -800 146022 480 0 FreeSans 1120 90 0 0 la_oenb[5]
port 503 nsew signal input
flabel metal2 s 340940 -800 341052 480 0 FreeSans 1120 90 0 0 la_oenb[60]
port 504 nsew signal input
flabel metal2 s 344486 -800 344598 480 0 FreeSans 1120 90 0 0 la_oenb[61]
port 505 nsew signal input
flabel metal2 s 348032 -800 348144 480 0 FreeSans 1120 90 0 0 la_oenb[62]
port 506 nsew signal input
flabel metal2 s 351578 -800 351690 480 0 FreeSans 1120 90 0 0 la_oenb[63]
port 507 nsew signal input
flabel metal2 s 355124 -800 355236 480 0 FreeSans 1120 90 0 0 la_oenb[64]
port 508 nsew signal input
flabel metal2 s 358670 -800 358782 480 0 FreeSans 1120 90 0 0 la_oenb[65]
port 509 nsew signal input
flabel metal2 s 362216 -800 362328 480 0 FreeSans 1120 90 0 0 la_oenb[66]
port 510 nsew signal input
flabel metal2 s 365762 -800 365874 480 0 FreeSans 1120 90 0 0 la_oenb[67]
port 511 nsew signal input
flabel metal2 s 369308 -800 369420 480 0 FreeSans 1120 90 0 0 la_oenb[68]
port 512 nsew signal input
flabel metal2 s 372854 -800 372966 480 0 FreeSans 1120 90 0 0 la_oenb[69]
port 513 nsew signal input
flabel metal2 s 149456 -800 149568 480 0 FreeSans 1120 90 0 0 la_oenb[6]
port 514 nsew signal input
flabel metal2 s 376400 -800 376512 480 0 FreeSans 1120 90 0 0 la_oenb[70]
port 515 nsew signal input
flabel metal2 s 379946 -800 380058 480 0 FreeSans 1120 90 0 0 la_oenb[71]
port 516 nsew signal input
flabel metal2 s 383492 -800 383604 480 0 FreeSans 1120 90 0 0 la_oenb[72]
port 517 nsew signal input
flabel metal2 s 387038 -800 387150 480 0 FreeSans 1120 90 0 0 la_oenb[73]
port 518 nsew signal input
flabel metal2 s 390584 -800 390696 480 0 FreeSans 1120 90 0 0 la_oenb[74]
port 519 nsew signal input
flabel metal2 s 394130 -800 394242 480 0 FreeSans 1120 90 0 0 la_oenb[75]
port 520 nsew signal input
flabel metal2 s 397676 -800 397788 480 0 FreeSans 1120 90 0 0 la_oenb[76]
port 521 nsew signal input
flabel metal2 s 401222 -800 401334 480 0 FreeSans 1120 90 0 0 la_oenb[77]
port 522 nsew signal input
flabel metal2 s 404768 -800 404880 480 0 FreeSans 1120 90 0 0 la_oenb[78]
port 523 nsew signal input
flabel metal2 s 408314 -800 408426 480 0 FreeSans 1120 90 0 0 la_oenb[79]
port 524 nsew signal input
flabel metal2 s 153002 -800 153114 480 0 FreeSans 1120 90 0 0 la_oenb[7]
port 525 nsew signal input
flabel metal2 s 411860 -800 411972 480 0 FreeSans 1120 90 0 0 la_oenb[80]
port 526 nsew signal input
flabel metal2 s 415406 -800 415518 480 0 FreeSans 1120 90 0 0 la_oenb[81]
port 527 nsew signal input
flabel metal2 s 418952 -800 419064 480 0 FreeSans 1120 90 0 0 la_oenb[82]
port 528 nsew signal input
flabel metal2 s 422498 -800 422610 480 0 FreeSans 1120 90 0 0 la_oenb[83]
port 529 nsew signal input
flabel metal2 s 426044 -800 426156 480 0 FreeSans 1120 90 0 0 la_oenb[84]
port 530 nsew signal input
flabel metal2 s 429590 -800 429702 480 0 FreeSans 1120 90 0 0 la_oenb[85]
port 531 nsew signal input
flabel metal2 s 433136 -800 433248 480 0 FreeSans 1120 90 0 0 la_oenb[86]
port 532 nsew signal input
flabel metal2 s 436682 -800 436794 480 0 FreeSans 1120 90 0 0 la_oenb[87]
port 533 nsew signal input
flabel metal2 s 440228 -800 440340 480 0 FreeSans 1120 90 0 0 la_oenb[88]
port 534 nsew signal input
flabel metal2 s 443774 -800 443886 480 0 FreeSans 1120 90 0 0 la_oenb[89]
port 535 nsew signal input
flabel metal2 s 156548 -800 156660 480 0 FreeSans 1120 90 0 0 la_oenb[8]
port 536 nsew signal input
flabel metal2 s 447320 -800 447432 480 0 FreeSans 1120 90 0 0 la_oenb[90]
port 537 nsew signal input
flabel metal2 s 450866 -800 450978 480 0 FreeSans 1120 90 0 0 la_oenb[91]
port 538 nsew signal input
flabel metal2 s 454412 -800 454524 480 0 FreeSans 1120 90 0 0 la_oenb[92]
port 539 nsew signal input
flabel metal2 s 457958 -800 458070 480 0 FreeSans 1120 90 0 0 la_oenb[93]
port 540 nsew signal input
flabel metal2 s 461504 -800 461616 480 0 FreeSans 1120 90 0 0 la_oenb[94]
port 541 nsew signal input
flabel metal2 s 465050 -800 465162 480 0 FreeSans 1120 90 0 0 la_oenb[95]
port 542 nsew signal input
flabel metal2 s 468596 -800 468708 480 0 FreeSans 1120 90 0 0 la_oenb[96]
port 543 nsew signal input
flabel metal2 s 472142 -800 472254 480 0 FreeSans 1120 90 0 0 la_oenb[97]
port 544 nsew signal input
flabel metal2 s 475688 -800 475800 480 0 FreeSans 1120 90 0 0 la_oenb[98]
port 545 nsew signal input
flabel metal2 s 479234 -800 479346 480 0 FreeSans 1120 90 0 0 la_oenb[99]
port 546 nsew signal input
flabel metal2 s 160094 -800 160206 480 0 FreeSans 1120 90 0 0 la_oenb[9]
port 547 nsew signal input
flabel metal2 s 579704 -800 579816 480 0 FreeSans 1120 90 0 0 user_clock2
port 548 nsew signal input
flabel metal2 s 580886 -800 580998 480 0 FreeSans 1120 90 0 0 user_irq[0]
port 549 nsew signal tristate
flabel metal2 s 582068 -800 582180 480 0 FreeSans 1120 90 0 0 user_irq[1]
port 550 nsew signal tristate
flabel metal2 s 583250 -800 583362 480 0 FreeSans 1120 90 0 0 user_irq[2]
port 551 nsew signal tristate
flabel metal3 s 582340 639784 584800 644584 0 FreeSans 1120 0 0 0 vccd1
port 552 nsew signal bidirectional
flabel metal3 s 582340 629784 584800 634584 0 FreeSans 1120 0 0 0 vccd1
port 553 nsew signal bidirectional
flabel metal3 s 0 643842 1660 648642 0 FreeSans 1120 0 0 0 vccd2
port 554 nsew signal bidirectional
flabel metal3 s 0 633842 1660 638642 0 FreeSans 1120 0 0 0 vccd2
port 555 nsew signal bidirectional
flabel metal3 s 582340 540562 584800 545362 0 FreeSans 1120 0 0 0 vdda1
port 556 nsew signal bidirectional
flabel metal3 s 582340 550562 584800 555362 0 FreeSans 1120 0 0 0 vdda1
port 557 nsew signal bidirectional
flabel metal3 s 582340 235230 584800 240030 0 FreeSans 1120 0 0 0 vdda1
port 558 nsew signal bidirectional
flabel metal3 s 582340 225230 584800 230030 0 FreeSans 1120 0 0 0 vdda1
port 559 nsew signal bidirectional
flabel metal3 s 0 204888 1660 209688 0 FreeSans 1120 0 0 0 vdda2
port 560 nsew signal bidirectional
flabel metal3 s 0 214888 1660 219688 0 FreeSans 1120 0 0 0 vdda2
port 561 nsew signal bidirectional
flabel metal3 s 520594 702340 525394 704800 0 FreeSans 1920 180 0 0 vssa1
port 562 nsew signal bidirectional
flabel metal3 s 510594 702340 515394 704800 0 FreeSans 1920 180 0 0 vssa1
port 563 nsew signal bidirectional
flabel metal3 s 582340 146830 584800 151630 0 FreeSans 1120 0 0 0 vssa1
port 564 nsew signal bidirectional
flabel metal3 s 582340 136830 584800 141630 0 FreeSans 1120 0 0 0 vssa1
port 565 nsew signal bidirectional
flabel metal3 s 0 559442 1660 564242 0 FreeSans 1120 0 0 0 vssa2
port 566 nsew signal bidirectional
flabel metal3 s 0 549442 1660 554242 0 FreeSans 1120 0 0 0 vssa2
port 567 nsew signal bidirectional
flabel metal3 s 0 172888 1660 177688 0 FreeSans 1120 0 0 0 vssd2
port 570 nsew signal bidirectional
flabel metal3 s 0 162888 1660 167688 0 FreeSans 1120 0 0 0 vssd2
port 571 nsew signal bidirectional
flabel metal2 s 524 -800 636 480 0 FreeSans 1120 90 0 0 wb_clk_i
port 572 nsew signal input
flabel metal2 s 1706 -800 1818 480 0 FreeSans 1120 90 0 0 wb_rst_i
port 573 nsew signal input
flabel metal2 s 2888 -800 3000 480 0 FreeSans 1120 90 0 0 wbs_ack_o
port 574 nsew signal tristate
flabel metal2 s 7616 -800 7728 480 0 FreeSans 1120 90 0 0 wbs_adr_i[0]
port 575 nsew signal input
flabel metal2 s 47804 -800 47916 480 0 FreeSans 1120 90 0 0 wbs_adr_i[10]
port 576 nsew signal input
flabel metal2 s 51350 -800 51462 480 0 FreeSans 1120 90 0 0 wbs_adr_i[11]
port 577 nsew signal input
flabel metal2 s 54896 -800 55008 480 0 FreeSans 1120 90 0 0 wbs_adr_i[12]
port 578 nsew signal input
flabel metal2 s 58442 -800 58554 480 0 FreeSans 1120 90 0 0 wbs_adr_i[13]
port 579 nsew signal input
flabel metal2 s 61988 -800 62100 480 0 FreeSans 1120 90 0 0 wbs_adr_i[14]
port 580 nsew signal input
flabel metal2 s 65534 -800 65646 480 0 FreeSans 1120 90 0 0 wbs_adr_i[15]
port 581 nsew signal input
flabel metal2 s 69080 -800 69192 480 0 FreeSans 1120 90 0 0 wbs_adr_i[16]
port 582 nsew signal input
flabel metal2 s 72626 -800 72738 480 0 FreeSans 1120 90 0 0 wbs_adr_i[17]
port 583 nsew signal input
flabel metal2 s 76172 -800 76284 480 0 FreeSans 1120 90 0 0 wbs_adr_i[18]
port 584 nsew signal input
flabel metal2 s 79718 -800 79830 480 0 FreeSans 1120 90 0 0 wbs_adr_i[19]
port 585 nsew signal input
flabel metal2 s 12344 -800 12456 480 0 FreeSans 1120 90 0 0 wbs_adr_i[1]
port 586 nsew signal input
flabel metal2 s 83264 -800 83376 480 0 FreeSans 1120 90 0 0 wbs_adr_i[20]
port 587 nsew signal input
flabel metal2 s 86810 -800 86922 480 0 FreeSans 1120 90 0 0 wbs_adr_i[21]
port 588 nsew signal input
flabel metal2 s 90356 -800 90468 480 0 FreeSans 1120 90 0 0 wbs_adr_i[22]
port 589 nsew signal input
flabel metal2 s 93902 -800 94014 480 0 FreeSans 1120 90 0 0 wbs_adr_i[23]
port 590 nsew signal input
flabel metal2 s 97448 -800 97560 480 0 FreeSans 1120 90 0 0 wbs_adr_i[24]
port 591 nsew signal input
flabel metal2 s 100994 -800 101106 480 0 FreeSans 1120 90 0 0 wbs_adr_i[25]
port 592 nsew signal input
flabel metal2 s 104540 -800 104652 480 0 FreeSans 1120 90 0 0 wbs_adr_i[26]
port 593 nsew signal input
flabel metal2 s 108086 -800 108198 480 0 FreeSans 1120 90 0 0 wbs_adr_i[27]
port 594 nsew signal input
flabel metal2 s 111632 -800 111744 480 0 FreeSans 1120 90 0 0 wbs_adr_i[28]
port 595 nsew signal input
flabel metal2 s 115178 -800 115290 480 0 FreeSans 1120 90 0 0 wbs_adr_i[29]
port 596 nsew signal input
flabel metal2 s 17072 -800 17184 480 0 FreeSans 1120 90 0 0 wbs_adr_i[2]
port 597 nsew signal input
flabel metal2 s 118724 -800 118836 480 0 FreeSans 1120 90 0 0 wbs_adr_i[30]
port 598 nsew signal input
flabel metal2 s 122270 -800 122382 480 0 FreeSans 1120 90 0 0 wbs_adr_i[31]
port 599 nsew signal input
flabel metal2 s 21800 -800 21912 480 0 FreeSans 1120 90 0 0 wbs_adr_i[3]
port 600 nsew signal input
flabel metal2 s 26528 -800 26640 480 0 FreeSans 1120 90 0 0 wbs_adr_i[4]
port 601 nsew signal input
flabel metal2 s 30074 -800 30186 480 0 FreeSans 1120 90 0 0 wbs_adr_i[5]
port 602 nsew signal input
flabel metal2 s 33620 -800 33732 480 0 FreeSans 1120 90 0 0 wbs_adr_i[6]
port 603 nsew signal input
flabel metal2 s 37166 -800 37278 480 0 FreeSans 1120 90 0 0 wbs_adr_i[7]
port 604 nsew signal input
flabel metal2 s 40712 -800 40824 480 0 FreeSans 1120 90 0 0 wbs_adr_i[8]
port 605 nsew signal input
flabel metal2 s 44258 -800 44370 480 0 FreeSans 1120 90 0 0 wbs_adr_i[9]
port 606 nsew signal input
flabel metal2 s 4070 -800 4182 480 0 FreeSans 1120 90 0 0 wbs_cyc_i
port 607 nsew signal input
flabel metal2 s 8798 -800 8910 480 0 FreeSans 1120 90 0 0 wbs_dat_i[0]
port 608 nsew signal input
flabel metal2 s 48986 -800 49098 480 0 FreeSans 1120 90 0 0 wbs_dat_i[10]
port 609 nsew signal input
flabel metal2 s 52532 -800 52644 480 0 FreeSans 1120 90 0 0 wbs_dat_i[11]
port 610 nsew signal input
flabel metal2 s 56078 -800 56190 480 0 FreeSans 1120 90 0 0 wbs_dat_i[12]
port 611 nsew signal input
flabel metal2 s 59624 -800 59736 480 0 FreeSans 1120 90 0 0 wbs_dat_i[13]
port 612 nsew signal input
flabel metal2 s 63170 -800 63282 480 0 FreeSans 1120 90 0 0 wbs_dat_i[14]
port 613 nsew signal input
flabel metal2 s 66716 -800 66828 480 0 FreeSans 1120 90 0 0 wbs_dat_i[15]
port 614 nsew signal input
flabel metal2 s 70262 -800 70374 480 0 FreeSans 1120 90 0 0 wbs_dat_i[16]
port 615 nsew signal input
flabel metal2 s 73808 -800 73920 480 0 FreeSans 1120 90 0 0 wbs_dat_i[17]
port 616 nsew signal input
flabel metal2 s 77354 -800 77466 480 0 FreeSans 1120 90 0 0 wbs_dat_i[18]
port 617 nsew signal input
flabel metal2 s 80900 -800 81012 480 0 FreeSans 1120 90 0 0 wbs_dat_i[19]
port 618 nsew signal input
flabel metal2 s 13526 -800 13638 480 0 FreeSans 1120 90 0 0 wbs_dat_i[1]
port 619 nsew signal input
flabel metal2 s 84446 -800 84558 480 0 FreeSans 1120 90 0 0 wbs_dat_i[20]
port 620 nsew signal input
flabel metal2 s 87992 -800 88104 480 0 FreeSans 1120 90 0 0 wbs_dat_i[21]
port 621 nsew signal input
flabel metal2 s 91538 -800 91650 480 0 FreeSans 1120 90 0 0 wbs_dat_i[22]
port 622 nsew signal input
flabel metal2 s 95084 -800 95196 480 0 FreeSans 1120 90 0 0 wbs_dat_i[23]
port 623 nsew signal input
flabel metal2 s 98630 -800 98742 480 0 FreeSans 1120 90 0 0 wbs_dat_i[24]
port 624 nsew signal input
flabel metal2 s 102176 -800 102288 480 0 FreeSans 1120 90 0 0 wbs_dat_i[25]
port 625 nsew signal input
flabel metal2 s 105722 -800 105834 480 0 FreeSans 1120 90 0 0 wbs_dat_i[26]
port 626 nsew signal input
flabel metal2 s 109268 -800 109380 480 0 FreeSans 1120 90 0 0 wbs_dat_i[27]
port 627 nsew signal input
flabel metal2 s 112814 -800 112926 480 0 FreeSans 1120 90 0 0 wbs_dat_i[28]
port 628 nsew signal input
flabel metal2 s 116360 -800 116472 480 0 FreeSans 1120 90 0 0 wbs_dat_i[29]
port 629 nsew signal input
flabel metal2 s 18254 -800 18366 480 0 FreeSans 1120 90 0 0 wbs_dat_i[2]
port 630 nsew signal input
flabel metal2 s 119906 -800 120018 480 0 FreeSans 1120 90 0 0 wbs_dat_i[30]
port 631 nsew signal input
flabel metal2 s 123452 -800 123564 480 0 FreeSans 1120 90 0 0 wbs_dat_i[31]
port 632 nsew signal input
flabel metal2 s 22982 -800 23094 480 0 FreeSans 1120 90 0 0 wbs_dat_i[3]
port 633 nsew signal input
flabel metal2 s 27710 -800 27822 480 0 FreeSans 1120 90 0 0 wbs_dat_i[4]
port 634 nsew signal input
flabel metal2 s 31256 -800 31368 480 0 FreeSans 1120 90 0 0 wbs_dat_i[5]
port 635 nsew signal input
flabel metal2 s 34802 -800 34914 480 0 FreeSans 1120 90 0 0 wbs_dat_i[6]
port 636 nsew signal input
flabel metal2 s 38348 -800 38460 480 0 FreeSans 1120 90 0 0 wbs_dat_i[7]
port 637 nsew signal input
flabel metal2 s 41894 -800 42006 480 0 FreeSans 1120 90 0 0 wbs_dat_i[8]
port 638 nsew signal input
flabel metal2 s 45440 -800 45552 480 0 FreeSans 1120 90 0 0 wbs_dat_i[9]
port 639 nsew signal input
flabel metal2 s 9980 -800 10092 480 0 FreeSans 1120 90 0 0 wbs_dat_o[0]
port 640 nsew signal tristate
flabel metal2 s 50168 -800 50280 480 0 FreeSans 1120 90 0 0 wbs_dat_o[10]
port 641 nsew signal tristate
flabel metal2 s 53714 -800 53826 480 0 FreeSans 1120 90 0 0 wbs_dat_o[11]
port 642 nsew signal tristate
flabel metal2 s 57260 -800 57372 480 0 FreeSans 1120 90 0 0 wbs_dat_o[12]
port 643 nsew signal tristate
flabel metal2 s 60806 -800 60918 480 0 FreeSans 1120 90 0 0 wbs_dat_o[13]
port 644 nsew signal tristate
flabel metal2 s 64352 -800 64464 480 0 FreeSans 1120 90 0 0 wbs_dat_o[14]
port 645 nsew signal tristate
flabel metal2 s 67898 -800 68010 480 0 FreeSans 1120 90 0 0 wbs_dat_o[15]
port 646 nsew signal tristate
flabel metal2 s 71444 -800 71556 480 0 FreeSans 1120 90 0 0 wbs_dat_o[16]
port 647 nsew signal tristate
flabel metal2 s 74990 -800 75102 480 0 FreeSans 1120 90 0 0 wbs_dat_o[17]
port 648 nsew signal tristate
flabel metal2 s 78536 -800 78648 480 0 FreeSans 1120 90 0 0 wbs_dat_o[18]
port 649 nsew signal tristate
flabel metal2 s 82082 -800 82194 480 0 FreeSans 1120 90 0 0 wbs_dat_o[19]
port 650 nsew signal tristate
flabel metal2 s 14708 -800 14820 480 0 FreeSans 1120 90 0 0 wbs_dat_o[1]
port 651 nsew signal tristate
flabel metal2 s 85628 -800 85740 480 0 FreeSans 1120 90 0 0 wbs_dat_o[20]
port 652 nsew signal tristate
flabel metal2 s 89174 -800 89286 480 0 FreeSans 1120 90 0 0 wbs_dat_o[21]
port 653 nsew signal tristate
flabel metal2 s 92720 -800 92832 480 0 FreeSans 1120 90 0 0 wbs_dat_o[22]
port 654 nsew signal tristate
flabel metal2 s 96266 -800 96378 480 0 FreeSans 1120 90 0 0 wbs_dat_o[23]
port 655 nsew signal tristate
flabel metal2 s 99812 -800 99924 480 0 FreeSans 1120 90 0 0 wbs_dat_o[24]
port 656 nsew signal tristate
flabel metal2 s 103358 -800 103470 480 0 FreeSans 1120 90 0 0 wbs_dat_o[25]
port 657 nsew signal tristate
flabel metal2 s 106904 -800 107016 480 0 FreeSans 1120 90 0 0 wbs_dat_o[26]
port 658 nsew signal tristate
flabel metal2 s 110450 -800 110562 480 0 FreeSans 1120 90 0 0 wbs_dat_o[27]
port 659 nsew signal tristate
flabel metal2 s 113996 -800 114108 480 0 FreeSans 1120 90 0 0 wbs_dat_o[28]
port 660 nsew signal tristate
flabel metal2 s 117542 -800 117654 480 0 FreeSans 1120 90 0 0 wbs_dat_o[29]
port 661 nsew signal tristate
flabel metal2 s 19436 -800 19548 480 0 FreeSans 1120 90 0 0 wbs_dat_o[2]
port 662 nsew signal tristate
flabel metal2 s 121088 -800 121200 480 0 FreeSans 1120 90 0 0 wbs_dat_o[30]
port 663 nsew signal tristate
flabel metal2 s 124634 -800 124746 480 0 FreeSans 1120 90 0 0 wbs_dat_o[31]
port 664 nsew signal tristate
flabel metal2 s 24164 -800 24276 480 0 FreeSans 1120 90 0 0 wbs_dat_o[3]
port 665 nsew signal tristate
flabel metal2 s 28892 -800 29004 480 0 FreeSans 1120 90 0 0 wbs_dat_o[4]
port 666 nsew signal tristate
flabel metal2 s 32438 -800 32550 480 0 FreeSans 1120 90 0 0 wbs_dat_o[5]
port 667 nsew signal tristate
flabel metal2 s 35984 -800 36096 480 0 FreeSans 1120 90 0 0 wbs_dat_o[6]
port 668 nsew signal tristate
flabel metal2 s 39530 -800 39642 480 0 FreeSans 1120 90 0 0 wbs_dat_o[7]
port 669 nsew signal tristate
flabel metal2 s 43076 -800 43188 480 0 FreeSans 1120 90 0 0 wbs_dat_o[8]
port 670 nsew signal tristate
flabel metal2 s 46622 -800 46734 480 0 FreeSans 1120 90 0 0 wbs_dat_o[9]
port 671 nsew signal tristate
flabel metal2 s 11162 -800 11274 480 0 FreeSans 1120 90 0 0 wbs_sel_i[0]
port 672 nsew signal input
flabel metal2 s 15890 -800 16002 480 0 FreeSans 1120 90 0 0 wbs_sel_i[1]
port 673 nsew signal input
flabel metal2 s 20618 -800 20730 480 0 FreeSans 1120 90 0 0 wbs_sel_i[2]
port 674 nsew signal input
flabel metal2 s 25346 -800 25458 480 0 FreeSans 1120 90 0 0 wbs_sel_i[3]
port 675 nsew signal input
flabel metal2 s 5252 -800 5364 480 0 FreeSans 1120 90 0 0 wbs_stb_i
port 676 nsew signal input
flabel metal2 s 6434 -800 6546 480 0 FreeSans 1120 90 0 0 wbs_we_i
port 677 nsew signal input
flabel metal3 s 582340 181430 584800 186230 0 FreeSans 1120 0 0 0 vssd1
port 569 nsew signal bidirectional
flabel metal3 s 582340 191430 584800 196230 0 FreeSans 1120 0 0 0 vssd1
port 568 nsew signal bidirectional
rlabel metal4 559206 641470 559206 641470 1 VDD
rlabel metal5 524812 682428 524812 682428 3 GND
rlabel metal5 165552 699664 165552 699664 7 Vn
rlabel metal5 217310 693970 217310 693970 7 Vp
rlabel metal3 68152 698908 68152 698908 7 CLK
rlabel metal3 465398 698900 465398 698900 7 Outp
rlabel metal3 413390 699678 413390 699678 7 Outn
rlabel metal3 438920 662050 438920 662050 7 L1
rlabel metal3 447318 662074 447318 662074 7 L2
flabel metal3 s 120194 702300 125194 704800 0 FreeSans 1920 180 0 0 io_analog[7]
port 44 nsew signal bidirectional
rlabel locali 107246 567078 107246 567078 7 GND
rlabel locali 107734 567078 107734 567078 7 GND
rlabel locali 101256 567116 101256 567116 7 GND
rlabel locali 101744 567116 101744 567116 7 GND
rlabel metal3 120172 691326 120172 691326 3 CLKBAR
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>
