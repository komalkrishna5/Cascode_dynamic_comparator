magic
tech sky130A
magscale 1 2
timestamp 1654340384
<< nwell >>
rect 415108 688720 415488 688888
rect 415108 686652 415228 688720
rect 569596 688682 569878 688684
rect 569596 688404 569920 688682
rect 569694 688330 569784 688404
rect 415108 686634 415410 686652
rect 415450 686636 415470 686640
rect 415108 686624 415488 686634
rect 415106 686340 415488 686624
rect 466974 686458 467294 686682
rect 70778 673802 71096 673962
rect 70788 673782 71096 673802
rect 70806 673776 71078 673782
rect 71044 673739 71078 673776
rect 122758 673528 123082 673738
rect 440058 591014 440376 591302
rect 448410 591030 448734 591294
rect 408706 587622 409044 587940
rect 408694 585520 408968 585840
<< pwell >>
rect 125134 694640 125776 694988
rect 73140 686438 73778 686980
rect 415534 688716 415722 688870
rect 415544 688590 415698 688716
rect 569316 688586 569542 688714
rect 569318 688294 569542 688586
rect 467352 686498 467522 686728
rect 70480 673296 70722 673462
rect 122548 673038 122704 673200
rect 440480 591110 440636 591312
rect 448836 591186 448968 591338
rect 406400 587394 406680 587556
rect 406440 585304 406674 585460
<< psubdiff >>
rect 125346 694758 125370 694852
rect 125578 694758 125602 694852
rect 415572 688744 415596 688792
rect 415678 688744 415702 688792
rect 569352 688490 569376 688548
rect 569474 688490 569498 688548
rect 73332 686672 73356 686780
rect 73570 686672 73594 686780
rect 467370 686592 467394 686640
rect 467476 686592 467500 686640
rect 70532 673316 70556 673364
rect 70682 673316 70706 673364
rect 122550 673072 122574 673118
rect 122670 673072 122694 673118
rect 448834 591232 448858 591280
rect 448952 591232 448976 591280
rect 440494 591184 440518 591232
rect 440604 591184 440628 591232
rect 406548 587500 406600 587524
rect 406548 587392 406600 587416
rect 421984 585556 422008 585642
rect 422150 585556 422174 585642
rect 406522 585420 406578 585444
rect 406522 585314 406578 585338
<< nsubdiff >>
rect 569646 688494 569670 688568
rect 569834 688494 569858 688568
rect 467044 686534 467068 686592
rect 467202 686534 467226 686592
rect 415174 686450 415198 686512
rect 415338 686450 415362 686512
rect 70824 673848 70848 673896
rect 70976 673848 71000 673896
rect 122842 673596 122866 673650
rect 123004 673596 123028 673650
rect 440104 591072 440128 591138
rect 440266 591072 440290 591138
rect 448478 591098 448502 591158
rect 448640 591098 448664 591158
rect 408830 587846 408894 587870
rect 408830 587678 408894 587702
rect 408794 585778 408858 585802
rect 408794 585596 408858 585620
<< psubdiffcont >>
rect 125370 694758 125578 694852
rect 415596 688744 415678 688792
rect 569376 688490 569474 688548
rect 73356 686672 73570 686780
rect 467394 686592 467476 686640
rect 70556 673316 70682 673364
rect 122574 673072 122670 673118
rect 448858 591232 448952 591280
rect 440518 591184 440604 591232
rect 406548 587416 406600 587500
rect 422008 585556 422150 585642
rect 406522 585338 406578 585420
<< nsubdiffcont >>
rect 569670 688494 569834 688568
rect 467068 686534 467202 686592
rect 415198 686450 415338 686512
rect 70848 673848 70976 673896
rect 122866 673596 123004 673650
rect 440128 591072 440266 591138
rect 448502 591098 448640 591158
rect 408830 587702 408894 587846
rect 408794 585620 408858 585778
<< locali >>
rect 119054 695204 119058 695352
rect 119054 694860 119226 695204
rect 119054 694852 125608 694860
rect 119054 694758 125370 694852
rect 125578 694758 125608 694852
rect 119054 694752 125608 694758
rect 467252 691416 467818 691454
rect 415410 691358 415468 691360
rect 415348 691316 415914 691358
rect 415348 691208 415392 691316
rect 415494 691208 415752 691316
rect 415854 691208 415914 691316
rect 415348 691076 415914 691208
rect 415348 690968 415392 691076
rect 415494 690968 415752 691076
rect 415854 690968 415914 691076
rect 467252 691308 467296 691416
rect 467398 691308 467656 691416
rect 467758 691308 467818 691416
rect 467252 691176 467818 691308
rect 467252 691068 467296 691176
rect 467398 691068 467656 691176
rect 467758 691068 467818 691176
rect 467252 691026 467818 691068
rect 569216 691416 569782 691454
rect 569216 691308 569260 691416
rect 569362 691308 569620 691416
rect 569722 691308 569782 691416
rect 569216 691176 569782 691308
rect 569216 691068 569260 691176
rect 569362 691068 569620 691176
rect 569722 691068 569782 691176
rect 569216 691028 569782 691068
rect 415348 690926 415914 690968
rect 415402 689342 415478 690926
rect 467318 690860 467482 691026
rect 415402 688666 415476 689342
rect 415580 688744 415596 688792
rect 415678 688744 415764 688792
rect 415408 688658 415474 688666
rect 412670 688608 414760 688612
rect 412670 688376 415068 688608
rect 415508 688595 415528 688670
rect 415728 688666 415764 688744
rect 467352 688664 467436 690860
rect 569394 690760 569728 691028
rect 569398 690550 569724 690760
rect 566276 689754 568936 689756
rect 566276 689750 568962 689754
rect 416130 688586 416872 688598
rect 412670 688212 413812 688376
rect 413996 688212 414212 688376
rect 414396 688212 415068 688376
rect 412670 687976 415068 688212
rect 412670 687812 413812 687976
rect 413996 687812 414212 687976
rect 414396 687812 415068 687976
rect 412670 687576 415068 687812
rect 67006 687402 67294 687430
rect 67006 687178 67028 687402
rect 67270 687178 67294 687402
rect 412670 687412 413812 687576
rect 413996 687412 414212 687576
rect 414396 687412 415068 687576
rect 67006 686784 67294 687178
rect 412670 687176 415068 687412
rect 412670 687012 413812 687176
rect 413996 687012 414212 687176
rect 414396 687012 415068 687176
rect 412670 686948 415068 687012
rect 416034 688376 416872 688586
rect 416034 688212 416278 688376
rect 416396 688212 416612 688376
rect 416796 688212 416872 688376
rect 416034 687976 416872 688212
rect 416034 687812 416278 687976
rect 416396 687812 416612 687976
rect 416796 687812 416872 687976
rect 416034 687576 416872 687812
rect 416034 687412 416278 687576
rect 416396 687412 416612 687576
rect 416796 687412 416872 687576
rect 416034 687176 416872 687412
rect 416034 687012 416278 687176
rect 416396 687012 416622 687176
rect 416806 687012 416872 687176
rect 412670 686942 414760 686948
rect 416034 686944 416872 687012
rect 465730 688376 466492 688608
rect 468130 688586 468872 688598
rect 465730 688212 465812 688376
rect 465996 688212 466212 688376
rect 466396 688212 466492 688376
rect 465730 687976 466492 688212
rect 465730 687812 465812 687976
rect 465996 687812 466212 687976
rect 466396 687812 466492 687976
rect 465730 687576 466492 687812
rect 465730 687412 465812 687576
rect 465996 687412 466212 687576
rect 466396 687412 466492 687576
rect 465730 687176 466492 687412
rect 465730 687012 465812 687176
rect 465996 687012 466212 687176
rect 466396 687012 466492 687176
rect 465730 686944 466492 687012
rect 468104 688376 468872 688586
rect 468104 688212 468212 688376
rect 468396 688212 468612 688376
rect 468796 688212 468872 688376
rect 468104 687976 468872 688212
rect 468104 687812 468212 687976
rect 468396 687812 468612 687976
rect 468796 687812 468872 687976
rect 468104 687576 468872 687812
rect 468104 687412 468212 687576
rect 468396 687412 468612 687576
rect 468796 687412 468872 687576
rect 468104 687176 468872 687412
rect 468104 687012 468212 687176
rect 468396 687012 468622 687176
rect 468806 687012 468872 687176
rect 468104 686944 468872 687012
rect 566276 688376 568976 689750
rect 569394 689304 569724 690550
rect 570186 689894 571476 689920
rect 570186 689592 571544 689894
rect 569546 689018 569606 689304
rect 570186 689284 571002 689592
rect 571242 689284 571544 689592
rect 570186 688992 571544 689284
rect 569360 688542 569376 688548
rect 566276 688212 568212 688376
rect 568396 688212 568612 688376
rect 568796 688212 568976 688376
rect 569316 688490 569376 688542
rect 569474 688490 569490 688548
rect 569316 688328 569366 688490
rect 569558 688285 569592 688835
rect 569696 688568 569786 688730
rect 570186 688684 571002 688992
rect 571242 688684 571544 688992
rect 569646 688494 569670 688568
rect 569834 688494 569850 688568
rect 569694 688330 569784 688494
rect 570186 688392 571544 688684
rect 566276 687976 568976 688212
rect 566276 687812 568212 687976
rect 568396 687812 568612 687976
rect 568796 687812 568976 687976
rect 566276 687576 568976 687812
rect 566276 687412 568212 687576
rect 568396 687412 568612 687576
rect 568796 687412 568976 687576
rect 566276 687176 568976 687412
rect 566276 687012 568212 687176
rect 568396 687012 568622 687176
rect 568806 687012 568976 687176
rect 416034 686936 416238 686944
rect 468104 686936 468238 686944
rect 67006 686780 73574 686784
rect 67006 686672 73356 686780
rect 73570 686672 73586 686780
rect 67006 686666 73574 686672
rect 415184 686512 415220 686680
rect 415494 686612 415532 686696
rect 415494 686562 415684 686612
rect 415182 686450 415198 686512
rect 415338 686450 415354 686512
rect 415184 686448 415220 686450
rect 415624 685910 415684 686562
rect 466992 686592 467028 686714
rect 466992 686534 467068 686592
rect 467202 686534 467218 686592
rect 467304 686184 467342 686724
rect 467540 686640 467576 686714
rect 467378 686592 467394 686640
rect 467476 686592 467576 686640
rect 415624 685558 415682 685910
rect 467304 685580 467344 686184
rect 415562 685516 416128 685558
rect 415562 685408 415606 685516
rect 415708 685408 415966 685516
rect 416068 685408 416128 685516
rect 415562 685276 416128 685408
rect 415562 685168 415606 685276
rect 415708 685168 415966 685276
rect 416068 685168 416128 685276
rect 415562 685126 416128 685168
rect 467146 685554 467380 685580
rect 467146 685512 467712 685554
rect 467146 685404 467190 685512
rect 467292 685404 467550 685512
rect 467652 685404 467712 685512
rect 566276 685506 568976 687012
rect 570186 688084 571002 688392
rect 571242 688084 571544 688392
rect 570186 687792 571544 688084
rect 570186 687484 571002 687792
rect 571242 687484 571544 687792
rect 570186 687192 571544 687484
rect 570186 686884 571002 687192
rect 571242 686884 571544 687192
rect 570186 686592 571544 686884
rect 566276 685486 568936 685506
rect 467146 685272 467712 685404
rect 467146 685164 467190 685272
rect 467292 685164 467550 685272
rect 467652 685164 467712 685272
rect 467146 685122 467712 685164
rect 569520 684432 569604 686400
rect 570186 686284 571002 686592
rect 571242 686284 571544 686592
rect 570186 685992 571544 686284
rect 570186 685684 571002 685992
rect 571242 685684 571544 685992
rect 570186 684684 571544 685684
rect 570818 684672 571544 684684
rect 569522 684204 569604 684432
rect 569518 683852 569604 684204
rect 569216 683816 569782 683852
rect 569216 683708 569260 683816
rect 569362 683708 569620 683816
rect 569722 683708 569782 683816
rect 569216 683576 569782 683708
rect 569216 683468 569260 683576
rect 569362 683468 569620 683576
rect 569722 683468 569782 683576
rect 569216 683434 569782 683468
rect 122524 674974 123090 675016
rect 70536 674932 71102 674974
rect 70536 674824 70580 674932
rect 70682 674824 70940 674932
rect 71042 674824 71102 674932
rect 70536 674692 71102 674824
rect 70536 674584 70580 674692
rect 70682 674584 70940 674692
rect 71042 674584 71102 674692
rect 122524 674866 122568 674974
rect 122670 674866 122928 674974
rect 123030 674866 123090 674974
rect 122524 674734 123090 674866
rect 122524 674626 122568 674734
rect 122670 674626 122928 674734
rect 123030 674626 123090 674734
rect 122524 674586 123090 674626
rect 70536 674544 71102 674584
rect 70718 673688 70784 674544
rect 70832 673848 70848 673896
rect 70976 673848 71078 673896
rect 122700 673848 122770 674586
rect 71044 673739 71078 673848
rect 70574 673364 70658 673426
rect 70540 673316 70556 673364
rect 70682 673316 70698 673364
rect 70574 673314 70658 673316
rect 70736 673170 70778 673522
rect 122696 673464 122770 673848
rect 122832 673596 122866 673650
rect 123004 673596 123062 673650
rect 123028 673478 123062 673596
rect 70678 672410 70798 673170
rect 122578 673118 122670 673178
rect 122558 673072 122574 673118
rect 122670 673072 122686 673118
rect 122720 673002 122762 673284
rect 122782 673260 122824 673270
rect 122668 672416 122786 673002
rect 70678 672374 70796 672410
rect 122514 672374 123080 672416
rect 70526 672332 71092 672374
rect 70526 672224 70570 672332
rect 70672 672224 70930 672332
rect 71032 672224 71092 672332
rect 70526 672092 71092 672224
rect 70526 671984 70570 672092
rect 70672 671984 70930 672092
rect 71032 671984 71092 672092
rect 122514 672266 122558 672374
rect 122660 672266 122918 672374
rect 123020 672266 123080 672374
rect 122514 672134 123080 672266
rect 122514 672026 122558 672134
rect 122660 672026 122918 672134
rect 123020 672026 123080 672134
rect 122514 671986 123080 672026
rect 70526 671944 71092 671984
rect 440208 593684 440774 593726
rect 440208 593576 440252 593684
rect 440354 593576 440612 593684
rect 440714 593576 440774 593684
rect 440208 593444 440774 593576
rect 440208 593336 440252 593444
rect 440354 593336 440612 593444
rect 440714 593336 440774 593444
rect 440208 593296 440774 593336
rect 448556 593716 449122 593758
rect 448556 593608 448600 593716
rect 448702 593608 448960 593716
rect 449062 593608 449122 593716
rect 448556 593476 449122 593608
rect 448556 593368 448600 593476
rect 448702 593368 448960 593476
rect 449062 593368 449122 593476
rect 448556 593328 449122 593368
rect 440364 592984 440462 593296
rect 448712 593004 448810 593328
rect 440364 592962 440464 592984
rect 437730 592374 438598 592380
rect 437730 592148 438850 592374
rect 437730 591984 437812 592148
rect 437996 591984 438212 592148
rect 438396 591984 438850 592148
rect 440366 592010 440464 592962
rect 442232 592244 443072 592420
rect 442232 592080 442412 592244
rect 442596 592080 442812 592244
rect 442996 592080 443072 592244
rect 437730 591748 438850 591984
rect 437730 591584 437812 591748
rect 437996 591584 438212 591748
rect 438396 591584 438850 591748
rect 437730 591348 438850 591584
rect 440384 591530 440420 592010
rect 442232 591938 443072 592080
rect 442214 591844 443072 591938
rect 442214 591680 442412 591844
rect 442596 591680 442812 591844
rect 442996 591680 443072 591844
rect 442214 591444 443072 591680
rect 437730 591184 437812 591348
rect 437996 591184 438212 591348
rect 438396 591184 438850 591348
rect 437730 590948 438850 591184
rect 440076 591150 440112 591348
rect 440076 591138 440290 591150
rect 440076 591078 440128 591138
rect 440080 591072 440128 591078
rect 440266 591072 440290 591138
rect 437730 590784 437812 590948
rect 437996 590784 438212 590948
rect 438396 590784 438850 590948
rect 437730 590716 438850 590784
rect 438466 590706 438850 590716
rect 440368 590258 440442 591374
rect 440622 591232 440660 591310
rect 440478 591184 440518 591232
rect 440604 591184 440660 591232
rect 442214 591280 442412 591444
rect 442596 591280 442812 591444
rect 442996 591280 443072 591444
rect 442214 591044 443072 591280
rect 442214 590950 442412 591044
rect 442232 590880 442412 590950
rect 442596 590880 442822 591044
rect 443006 590880 443072 591044
rect 442232 590812 443072 590880
rect 446130 592374 446998 592380
rect 446130 592148 447250 592374
rect 446130 591984 446212 592148
rect 446396 591984 446612 592148
rect 446796 591984 447250 592148
rect 446130 591748 447250 591984
rect 448710 591922 448810 593004
rect 450694 592244 451472 592420
rect 450694 592080 450812 592244
rect 450996 592080 451212 592244
rect 451396 592080 451472 592244
rect 446130 591584 446212 591748
rect 446396 591584 446612 591748
rect 446796 591584 447250 591748
rect 446130 591348 447250 591584
rect 448736 591552 448774 591922
rect 450694 591844 451472 592080
rect 450694 591680 450812 591844
rect 450996 591680 451212 591844
rect 451396 591680 451472 591844
rect 450694 591444 451472 591680
rect 446130 591184 446212 591348
rect 446396 591184 446612 591348
rect 446796 591184 447250 591348
rect 446130 590948 447250 591184
rect 448430 591166 448466 591352
rect 448738 591342 448786 591396
rect 448430 591158 448662 591166
rect 448430 591098 448502 591158
rect 448640 591098 448662 591158
rect 442232 590804 442438 590812
rect 446130 590784 446212 590948
rect 446396 590784 446612 590948
rect 446796 590784 447250 590948
rect 446130 590716 447250 590784
rect 446866 590706 447250 590716
rect 448738 591002 448784 591342
rect 448974 591282 449014 591332
rect 448842 591232 448858 591280
rect 448952 591232 449014 591282
rect 450694 591280 450812 591444
rect 450996 591280 451212 591444
rect 451396 591280 451472 591444
rect 450694 591044 451472 591280
rect 448738 590332 448786 591002
rect 450694 590880 450812 591044
rect 450996 590880 451222 591044
rect 451406 590880 451472 591044
rect 450694 590812 451472 590880
rect 450694 590804 450838 590812
rect 440368 590254 440452 590258
rect 448696 590254 448814 590332
rect 440216 590212 440782 590254
rect 440216 590104 440260 590212
rect 440362 590104 440620 590212
rect 440722 590104 440782 590212
rect 440216 589972 440782 590104
rect 440216 589864 440260 589972
rect 440362 589864 440620 589972
rect 440722 589864 440782 589972
rect 440216 589824 440782 589864
rect 448544 590212 449110 590254
rect 448544 590104 448588 590212
rect 448690 590104 448948 590212
rect 449050 590104 449110 590212
rect 448544 589972 449110 590104
rect 448544 589864 448588 589972
rect 448690 589864 448948 589972
rect 449050 589864 449110 589972
rect 448544 589824 449110 589864
rect 405258 588544 410482 588850
rect 405258 588304 405560 588544
rect 405868 588304 406160 588544
rect 406468 588304 406760 588544
rect 407068 588304 407360 588544
rect 407668 588304 407960 588544
rect 408268 588304 408560 588544
rect 408868 588304 409160 588544
rect 409468 588304 410482 588544
rect 405258 588056 410482 588304
rect 408632 587882 408898 587922
rect 408830 587846 408894 587882
rect 404984 587696 405238 587706
rect 404984 587640 405006 587696
rect 405086 587640 405126 587696
rect 405206 587640 405238 587696
rect 408830 587686 408894 587702
rect 409968 587696 410212 587706
rect 409968 587646 409990 587696
rect 409966 587640 409990 587646
rect 410070 587640 410110 587696
rect 410190 587640 410212 587696
rect 404984 587634 405238 587640
rect 404984 587632 405336 587634
rect 404984 587614 406572 587632
rect 408624 587620 409758 587640
rect 409966 587620 410212 587640
rect 404984 587612 406634 587614
rect 404984 587596 406676 587612
rect 404984 587540 405006 587596
rect 405086 587540 405126 587596
rect 405206 587574 406676 587596
rect 408624 587596 410212 587620
rect 405206 587572 406634 587574
rect 405206 587556 406572 587572
rect 408624 587566 409990 587596
rect 405206 587554 405336 587556
rect 405206 587540 405238 587554
rect 404984 587510 405238 587540
rect 408624 587536 409758 587566
rect 409968 587540 409990 587566
rect 410070 587540 410110 587596
rect 410190 587540 410212 587596
rect 406548 587500 406600 587516
rect 409968 587510 410212 587540
rect 406600 587416 406712 587480
rect 406548 587400 406600 587416
rect 405234 587030 410098 587154
rect 405234 586866 405398 587030
rect 405592 586866 405798 587030
rect 405992 586866 406198 587030
rect 406392 586866 406598 587030
rect 406792 586866 406998 587030
rect 407192 586866 407398 587030
rect 407592 586866 407798 587030
rect 407992 586866 408198 587030
rect 408392 586866 408598 587030
rect 408792 586866 408998 587030
rect 409192 586866 409398 587030
rect 409592 586866 409798 587030
rect 409992 586866 410098 587030
rect 405234 586790 410098 586866
rect 405234 586626 405398 586790
rect 405592 586626 405798 586790
rect 405992 586626 406198 586790
rect 406392 586626 406598 586790
rect 406792 586626 406998 586790
rect 407192 586626 407398 586790
rect 407592 586626 407798 586790
rect 407992 586626 408198 586790
rect 408392 586626 408598 586790
rect 408792 586626 408998 586790
rect 409192 586626 409398 586790
rect 409592 586626 409798 586790
rect 409992 586626 410098 586790
rect 405234 586572 410098 586626
rect 405242 586562 410086 586572
rect 405396 586344 410074 586454
rect 405396 586104 405560 586344
rect 405868 586104 406160 586344
rect 406468 586104 406760 586344
rect 407068 586104 407360 586344
rect 407668 586104 407960 586344
rect 408268 586104 408560 586344
rect 408868 586104 409160 586344
rect 409468 586104 410074 586344
rect 405396 585978 410074 586104
rect 408640 585782 408858 585818
rect 408794 585778 408858 585782
rect 404984 585596 405258 585606
rect 408794 585604 408858 585620
rect 404984 585540 405006 585596
rect 405086 585540 405126 585596
rect 405206 585540 405258 585596
rect 409976 585596 410220 585606
rect 404984 585516 405258 585540
rect 408616 585544 408650 585584
rect 409976 585546 409998 585596
rect 409814 585544 409998 585546
rect 408616 585540 409998 585544
rect 410078 585540 410118 585596
rect 410198 585540 410220 585596
rect 421924 585556 422008 585642
rect 422150 585556 422166 585642
rect 404984 585512 406616 585516
rect 404984 585496 406668 585512
rect 404984 585440 405006 585496
rect 405086 585440 405126 585496
rect 405206 585470 406668 585496
rect 408616 585496 410220 585540
rect 405206 585440 405258 585470
rect 408616 585444 409998 585496
rect 404984 585410 405258 585440
rect 409976 585440 409998 585444
rect 410078 585440 410118 585496
rect 410198 585440 410220 585496
rect 406522 585420 406578 585436
rect 406578 585338 406692 585418
rect 409976 585410 410220 585440
rect 406522 585322 406578 585338
rect 405242 585030 410086 585078
rect 405242 584866 405398 585030
rect 405592 584866 405798 585030
rect 405992 584866 406198 585030
rect 406392 584866 406598 585030
rect 406792 584866 406998 585030
rect 407192 584866 407398 585030
rect 407592 584866 407798 585030
rect 407992 584866 408198 585030
rect 408392 584866 408598 585030
rect 408792 584866 408998 585030
rect 409192 584866 409398 585030
rect 409592 584866 409798 585030
rect 409992 584866 410086 585030
rect 405242 584790 410086 584866
rect 405242 584626 405398 584790
rect 405592 584626 405798 584790
rect 405992 584626 406198 584790
rect 406392 584626 406598 584790
rect 406792 584626 406998 584790
rect 407192 584626 407398 584790
rect 407592 584626 407798 584790
rect 407992 584626 408198 584790
rect 408392 584626 408598 584790
rect 408792 584626 408998 584790
rect 409192 584626 409398 584790
rect 409592 584626 409798 584790
rect 409992 584626 410086 584790
rect 405242 584562 410086 584626
<< viali >>
rect 119058 695204 119246 695372
rect 119380 695200 119414 695412
rect 125571 695233 125605 695335
rect 415392 691208 415494 691316
rect 415752 691208 415854 691316
rect 415392 690968 415494 691076
rect 415752 690968 415854 691076
rect 467296 691308 467398 691416
rect 467656 691308 467758 691416
rect 467296 691068 467398 691176
rect 467656 691068 467758 691176
rect 569260 691308 569362 691416
rect 569620 691308 569722 691416
rect 569260 691068 569362 691176
rect 569620 691068 569722 691176
rect 413812 688212 413996 688376
rect 414212 688212 414396 688376
rect 413812 687812 413996 687976
rect 414212 687812 414396 687976
rect 67028 687178 67270 687402
rect 413812 687412 413996 687576
rect 414212 687412 414396 687576
rect 67401 687251 67435 687353
rect 73573 687233 73607 687335
rect 413812 687012 413996 687176
rect 414212 687012 414396 687176
rect 416278 688212 416396 688376
rect 416612 688212 416796 688376
rect 416278 687812 416396 687976
rect 416612 687812 416796 687976
rect 416278 687412 416396 687576
rect 416612 687412 416796 687576
rect 416278 687012 416396 687176
rect 416622 687012 416806 687176
rect 465812 688212 465996 688376
rect 466212 688212 466396 688376
rect 465812 687812 465996 687976
rect 466212 687812 466396 687976
rect 465812 687412 465996 687576
rect 466212 687412 466396 687576
rect 465812 687012 465996 687176
rect 466212 687012 466396 687176
rect 468212 688212 468396 688376
rect 468612 688212 468796 688376
rect 468212 687812 468396 687976
rect 468612 687812 468796 687976
rect 468212 687412 468396 687576
rect 468612 687412 468796 687576
rect 468212 687012 468396 687176
rect 468622 687012 468806 687176
rect 571002 689284 571242 689592
rect 568212 688212 568396 688376
rect 568612 688212 568796 688376
rect 571002 688684 571242 688992
rect 568212 687812 568396 687976
rect 568612 687812 568796 687976
rect 568212 687412 568396 687576
rect 568612 687412 568796 687576
rect 568212 687012 568396 687176
rect 568622 687012 568806 687176
rect 415606 685408 415708 685516
rect 415966 685408 416068 685516
rect 415606 685168 415708 685276
rect 415966 685168 416068 685276
rect 467190 685404 467292 685512
rect 467550 685404 467652 685512
rect 571002 688084 571242 688392
rect 571002 687484 571242 687792
rect 571002 686884 571242 687192
rect 467190 685164 467292 685272
rect 467550 685164 467652 685272
rect 571002 686284 571242 686592
rect 571002 685684 571242 685992
rect 569260 683708 569362 683816
rect 569620 683708 569722 683816
rect 569260 683468 569362 683576
rect 569620 683468 569722 683576
rect 70580 674824 70682 674932
rect 70940 674824 71042 674932
rect 70580 674584 70682 674692
rect 70940 674584 71042 674692
rect 122568 674866 122670 674974
rect 122928 674866 123030 674974
rect 122568 674626 122670 674734
rect 122928 674626 123030 674734
rect 70570 672224 70672 672332
rect 70930 672224 71032 672332
rect 70570 671984 70672 672092
rect 70930 671984 71032 672092
rect 122558 672266 122660 672374
rect 122918 672266 123020 672374
rect 122558 672026 122660 672134
rect 122918 672026 123020 672134
rect 440252 593576 440354 593684
rect 440612 593576 440714 593684
rect 440252 593336 440354 593444
rect 440612 593336 440714 593444
rect 448600 593608 448702 593716
rect 448960 593608 449062 593716
rect 448600 593368 448702 593476
rect 448960 593368 449062 593476
rect 437812 591984 437996 592148
rect 438212 591984 438396 592148
rect 442412 592080 442596 592244
rect 442812 592080 442996 592244
rect 437812 591584 437996 591748
rect 438212 591584 438396 591748
rect 442412 591680 442596 591844
rect 442812 591680 442996 591844
rect 437812 591184 437996 591348
rect 438212 591184 438396 591348
rect 437812 590784 437996 590948
rect 438212 590784 438396 590948
rect 442412 591280 442596 591444
rect 442812 591280 442996 591444
rect 442412 590880 442596 591044
rect 442822 590880 443006 591044
rect 446212 591984 446396 592148
rect 446612 591984 446796 592148
rect 450812 592080 450996 592244
rect 451212 592080 451396 592244
rect 446212 591584 446396 591748
rect 446612 591584 446796 591748
rect 450812 591680 450996 591844
rect 451212 591680 451396 591844
rect 446212 591184 446396 591348
rect 446612 591184 446796 591348
rect 446212 590784 446396 590948
rect 446612 590784 446796 590948
rect 450812 591280 450996 591444
rect 451212 591280 451396 591444
rect 450812 590880 450996 591044
rect 451222 590880 451406 591044
rect 440260 590104 440362 590212
rect 440620 590104 440722 590212
rect 440260 589864 440362 589972
rect 440620 589864 440722 589972
rect 448588 590104 448690 590212
rect 448948 590104 449050 590212
rect 448588 589864 448690 589972
rect 448948 589864 449050 589972
rect 405560 588304 405868 588544
rect 406160 588304 406468 588544
rect 406760 588304 407068 588544
rect 407360 588304 407668 588544
rect 407960 588304 408268 588544
rect 408560 588304 408868 588544
rect 409160 588304 409468 588544
rect 405006 587640 405086 587696
rect 405126 587640 405206 587696
rect 409990 587640 410070 587696
rect 410110 587640 410190 587696
rect 405006 587540 405086 587596
rect 405126 587540 405206 587596
rect 409990 587540 410070 587596
rect 410110 587540 410190 587596
rect 405398 586866 405592 587030
rect 405798 586866 405992 587030
rect 406198 586866 406392 587030
rect 406598 586866 406792 587030
rect 406998 586866 407192 587030
rect 407398 586866 407592 587030
rect 407798 586866 407992 587030
rect 408198 586866 408392 587030
rect 408598 586866 408792 587030
rect 408998 586866 409192 587030
rect 409398 586866 409592 587030
rect 409798 586866 409992 587030
rect 405398 586626 405592 586790
rect 405798 586626 405992 586790
rect 406198 586626 406392 586790
rect 406598 586626 406792 586790
rect 406998 586626 407192 586790
rect 407398 586626 407592 586790
rect 407798 586626 407992 586790
rect 408198 586626 408392 586790
rect 408598 586626 408792 586790
rect 408998 586626 409192 586790
rect 409398 586626 409592 586790
rect 409798 586626 409992 586790
rect 405560 586104 405868 586344
rect 406160 586104 406468 586344
rect 406760 586104 407068 586344
rect 407360 586104 407668 586344
rect 407960 586104 408268 586344
rect 408560 586104 408868 586344
rect 409160 586104 409468 586344
rect 405006 585540 405086 585596
rect 405126 585540 405206 585596
rect 409998 585540 410078 585596
rect 410118 585540 410198 585596
rect 405006 585440 405086 585496
rect 405126 585440 405206 585496
rect 409998 585440 410078 585496
rect 410118 585440 410198 585496
rect 405398 584866 405592 585030
rect 405798 584866 405992 585030
rect 406198 584866 406392 585030
rect 406598 584866 406792 585030
rect 406998 584866 407192 585030
rect 407398 584866 407592 585030
rect 407798 584866 407992 585030
rect 408198 584866 408392 585030
rect 408598 584866 408792 585030
rect 408998 584866 409192 585030
rect 409398 584866 409592 585030
rect 409798 584866 409992 585030
rect 405398 584626 405592 584790
rect 405798 584626 405992 584790
rect 406198 584626 406392 584790
rect 406598 584626 406792 584790
rect 406998 584626 407192 584790
rect 407398 584626 407592 584790
rect 407798 584626 407992 584790
rect 408198 584626 408392 584790
rect 408598 584626 408792 584790
rect 408998 584626 409192 584790
rect 409398 584626 409592 584790
rect 409798 584626 409992 584790
<< metal1 >>
rect 118982 695430 119314 695452
rect 119474 695442 119988 695450
rect 120218 695446 124754 696194
rect 120218 695442 120660 695446
rect 118982 695156 119008 695430
rect 119292 695412 119428 695430
rect 119292 695200 119380 695412
rect 119414 695200 119428 695412
rect 119292 695186 119428 695200
rect 119292 695156 119314 695186
rect 119474 695160 120660 695442
rect 119474 695158 119988 695160
rect 118982 695134 119314 695156
rect 120218 694918 120660 695160
rect 121252 694918 121760 695446
rect 122352 694918 122860 695446
rect 123452 694918 123960 695446
rect 124552 695442 124754 695446
rect 126154 695464 126622 695526
rect 124552 695160 125518 695442
rect 125558 695416 125884 695418
rect 126154 695416 126230 695464
rect 125558 695335 126230 695416
rect 125558 695233 125571 695335
rect 125605 695233 126230 695335
rect 125558 695174 126230 695233
rect 125558 695172 125884 695174
rect 124552 694918 124754 695160
rect 124980 695152 125518 695160
rect 126154 695110 126230 695174
rect 126562 695110 126622 695464
rect 126154 695056 126622 695110
rect 120218 694338 124754 694918
rect 467252 691416 467818 691454
rect 415348 691316 415914 691358
rect 415348 691208 415392 691316
rect 415494 691208 415752 691316
rect 415854 691208 415914 691316
rect 415348 691076 415914 691208
rect 415348 690968 415392 691076
rect 415494 690968 415752 691076
rect 415854 690968 415914 691076
rect 467252 691308 467296 691416
rect 467398 691308 467656 691416
rect 467758 691308 467818 691416
rect 467252 691176 467818 691308
rect 467252 691068 467296 691176
rect 467398 691068 467656 691176
rect 467758 691068 467818 691176
rect 467252 691026 467818 691068
rect 569216 691416 569782 691454
rect 569216 691308 569260 691416
rect 569362 691308 569620 691416
rect 569722 691308 569782 691416
rect 569216 691176 569782 691308
rect 569216 691068 569260 691176
rect 569362 691068 569620 691176
rect 569722 691068 569782 691176
rect 569216 691028 569782 691068
rect 415348 690926 415914 690968
rect 570922 689592 571352 689764
rect 570922 689284 571002 689592
rect 571242 689284 571352 689592
rect 569882 689070 570312 689072
rect 570922 689070 571352 689284
rect 568938 689064 569332 689066
rect 568122 688696 569332 689064
rect 569882 689018 571436 689070
rect 569884 688992 571436 689018
rect 569884 688696 571002 688992
rect 413726 688376 415224 688616
rect 413726 688212 413812 688376
rect 413996 688212 414212 688376
rect 414396 688212 415224 688376
rect 66982 687430 67314 687452
rect 68218 687446 72754 688194
rect 413726 687976 415224 688212
rect 413726 687812 413812 687976
rect 413996 687812 414212 687976
rect 414396 687812 415224 687976
rect 413726 687576 415224 687812
rect 74154 687464 74622 687526
rect 73002 687450 73512 687454
rect 67374 687430 67448 687432
rect 66982 687156 67008 687430
rect 67292 687353 67448 687430
rect 68218 687384 68660 687446
rect 67874 687382 68660 687384
rect 67292 687251 67401 687353
rect 67435 687251 67448 687353
rect 67292 687186 67448 687251
rect 67498 687232 68660 687382
rect 67874 687230 68660 687232
rect 67292 687156 67314 687186
rect 66982 687134 67314 687156
rect 68218 686918 68660 687230
rect 69252 686918 69760 687446
rect 70352 686918 70860 687446
rect 71452 686918 71960 687446
rect 72552 687442 72754 687446
rect 72988 687442 73512 687450
rect 72552 687160 73512 687442
rect 74154 687416 74230 687464
rect 73566 687335 74230 687416
rect 73566 687233 73573 687335
rect 73607 687233 74230 687335
rect 73566 687174 74230 687233
rect 72552 686918 72754 687160
rect 72988 687158 73512 687160
rect 73002 687156 73512 687158
rect 74154 687110 74230 687174
rect 74562 687110 74622 687464
rect 74154 687056 74622 687110
rect 413726 687412 413812 687576
rect 413996 687412 414212 687576
rect 414396 687412 415224 687576
rect 413726 687176 415224 687412
rect 413726 687012 413812 687176
rect 413996 687012 414212 687176
rect 414396 687012 415224 687176
rect 413726 686942 415224 687012
rect 415772 688376 416876 688694
rect 467560 688624 467948 688632
rect 465760 688608 467008 688616
rect 415772 688212 416278 688376
rect 416396 688212 416612 688376
rect 416796 688212 416876 688376
rect 415772 687976 416876 688212
rect 415772 687812 416278 687976
rect 416396 687812 416612 687976
rect 416796 687812 416876 687976
rect 415772 687576 416876 687812
rect 415772 687412 416278 687576
rect 416396 687412 416612 687576
rect 416796 687412 416876 687576
rect 415772 687176 416876 687412
rect 415772 687012 416278 687176
rect 416396 687012 416622 687176
rect 416806 687012 416876 687176
rect 68218 686338 72754 686918
rect 415698 686666 415765 686784
rect 415772 686662 416876 687012
rect 465730 688376 467008 688608
rect 465730 688212 465812 688376
rect 465996 688212 466212 688376
rect 466396 688212 467008 688376
rect 465730 687976 467008 688212
rect 465730 687812 465812 687976
rect 465996 687812 466212 687976
rect 466396 687812 467008 687976
rect 465730 687576 467008 687812
rect 465730 687412 465812 687576
rect 465996 687412 466212 687576
rect 466396 687412 467008 687576
rect 465730 687176 467008 687412
rect 465730 687012 465812 687176
rect 465996 687012 466212 687176
rect 466396 687012 467008 687176
rect 465730 686944 467008 687012
rect 467560 688598 468828 688624
rect 467560 688376 468866 688598
rect 568122 688420 569218 688696
rect 569960 688684 571002 688696
rect 571242 688684 571436 688992
rect 568122 688410 569366 688420
rect 467560 688212 468212 688376
rect 468396 688212 468612 688376
rect 468796 688212 468866 688376
rect 467560 687976 468866 688212
rect 467560 687812 468212 687976
rect 468396 687812 468612 687976
rect 468796 687812 468866 687976
rect 467560 687576 468866 687812
rect 467560 687412 468212 687576
rect 468396 687412 468612 687576
rect 468796 687412 468866 687576
rect 467560 687176 468866 687412
rect 467560 687012 468212 687176
rect 468396 687012 468622 687176
rect 468806 687012 468866 687176
rect 467560 686956 468866 687012
rect 467560 686950 467948 686956
rect 468130 686944 468866 686956
rect 568128 688376 569366 688410
rect 569960 688392 571436 688684
rect 569960 688390 571002 688392
rect 568128 688212 568212 688376
rect 568396 688212 568612 688376
rect 568796 688212 569366 688376
rect 568128 687976 569366 688212
rect 568128 687812 568212 687976
rect 568396 687812 568612 687976
rect 568796 687812 569366 687976
rect 568128 687576 569366 687812
rect 568128 687412 568212 687576
rect 568396 687412 568612 687576
rect 568796 687412 569366 687576
rect 568128 687176 569366 687412
rect 568128 687012 568212 687176
rect 568396 687012 568622 687176
rect 568806 687012 569366 687176
rect 465760 686942 467008 686944
rect 568128 686370 569366 687012
rect 569880 688084 571002 688390
rect 571242 688390 571436 688392
rect 571242 688084 571438 688390
rect 569880 687792 571438 688084
rect 569880 687484 571002 687792
rect 571242 687484 571438 687792
rect 569880 687192 571438 687484
rect 569880 686884 571002 687192
rect 571242 686884 571438 687192
rect 569880 686592 571438 686884
rect 569880 686324 571002 686592
rect 570922 686284 571002 686324
rect 571242 686324 571438 686592
rect 571242 686284 571352 686324
rect 570922 685992 571352 686284
rect 570922 685684 571002 685992
rect 571242 685684 571352 685992
rect 415562 685516 416128 685558
rect 415562 685408 415606 685516
rect 415708 685408 415966 685516
rect 416068 685408 416128 685516
rect 415562 685276 416128 685408
rect 415562 685168 415606 685276
rect 415708 685168 415966 685276
rect 416068 685168 416128 685276
rect 415562 685126 416128 685168
rect 467146 685554 467272 685580
rect 467146 685512 467712 685554
rect 467146 685404 467190 685512
rect 467292 685404 467550 685512
rect 467652 685404 467712 685512
rect 467146 685272 467712 685404
rect 467146 685164 467190 685272
rect 467292 685164 467550 685272
rect 467652 685164 467712 685272
rect 467146 685122 467712 685164
rect 570922 685072 571352 685684
rect 569216 683816 569782 683852
rect 569216 683708 569260 683816
rect 569362 683708 569620 683816
rect 569722 683708 569782 683816
rect 569216 683576 569782 683708
rect 569216 683468 569260 683576
rect 569362 683468 569620 683576
rect 569722 683468 569782 683576
rect 569216 683434 569782 683468
rect 122524 674974 123090 675016
rect 70536 674932 71102 674974
rect 70536 674824 70580 674932
rect 70682 674824 70940 674932
rect 71042 674824 71102 674932
rect 70536 674692 71102 674824
rect 70536 674584 70580 674692
rect 70682 674584 70940 674692
rect 71042 674584 71102 674692
rect 122524 674866 122568 674974
rect 122670 674866 122928 674974
rect 123030 674866 123090 674974
rect 122524 674734 123090 674866
rect 122524 674626 122568 674734
rect 122670 674626 122928 674734
rect 123030 674626 123090 674734
rect 122524 674586 123090 674626
rect 70536 674544 71102 674584
rect 69934 673768 70382 673770
rect 69934 673732 70482 673768
rect 69934 673458 70008 673732
rect 70292 673724 70482 673732
rect 71292 673756 71760 673818
rect 70292 673458 70560 673724
rect 71292 673708 71368 673756
rect 71038 673466 71368 673708
rect 69934 673400 70560 673458
rect 71292 673402 71368 673466
rect 71700 673402 71760 673756
rect 69934 673398 70482 673400
rect 71292 673348 71760 673402
rect 121734 673518 122168 673532
rect 123226 673524 123694 673526
rect 121734 673516 122434 673518
rect 121734 673504 122466 673516
rect 121734 673498 122476 673504
rect 122526 673498 122548 673504
rect 121734 673494 122548 673498
rect 121734 673220 121808 673494
rect 122092 673220 122548 673494
rect 123082 673464 123694 673524
rect 123082 673416 123302 673464
rect 123020 673260 123302 673416
rect 121734 673160 122548 673220
rect 122058 673150 122548 673160
rect 123082 673150 123302 673260
rect 122058 673148 122298 673150
rect 122398 673148 122548 673150
rect 123226 673110 123302 673150
rect 123634 673110 123694 673464
rect 123226 673056 123694 673110
rect 122514 672374 123080 672416
rect 70526 672332 71092 672374
rect 70526 672224 70570 672332
rect 70672 672224 70930 672332
rect 71032 672224 71092 672332
rect 70526 672092 71092 672224
rect 70526 671984 70570 672092
rect 70672 671984 70930 672092
rect 71032 671984 71092 672092
rect 122514 672266 122558 672374
rect 122660 672266 122918 672374
rect 123020 672266 123080 672374
rect 122514 672134 123080 672266
rect 122514 672026 122558 672134
rect 122660 672026 122918 672134
rect 123020 672026 123080 672134
rect 122514 671986 123080 672026
rect 70526 671944 71092 671984
rect 440208 593684 440774 593726
rect 440208 593576 440252 593684
rect 440354 593576 440612 593684
rect 440714 593576 440774 593684
rect 440208 593444 440774 593576
rect 440208 593336 440252 593444
rect 440354 593336 440612 593444
rect 440714 593336 440774 593444
rect 440208 593296 440774 593336
rect 448556 593716 449122 593758
rect 448556 593608 448600 593716
rect 448702 593608 448960 593716
rect 449062 593608 449122 593716
rect 448556 593476 449122 593608
rect 448556 593368 448600 593476
rect 448702 593368 448960 593476
rect 449062 593368 449122 593476
rect 448556 593328 449122 593368
rect 442330 592416 443066 592420
rect 450730 592416 451466 592420
rect 437730 592148 440102 592380
rect 437730 591984 437812 592148
rect 437996 591984 438212 592148
rect 438396 591984 440102 592148
rect 437730 591748 440102 591984
rect 437730 591584 437812 591748
rect 437996 591584 438212 591748
rect 438396 591584 440102 591748
rect 437730 591348 440102 591584
rect 437730 591184 437812 591348
rect 437996 591184 438212 591348
rect 438396 591184 440102 591348
rect 437730 590948 440102 591184
rect 437730 590784 437812 590948
rect 437996 590784 438212 590948
rect 438396 590784 440102 590948
rect 437730 590716 440102 590784
rect 440650 592244 443196 592416
rect 440650 592080 442412 592244
rect 442596 592080 442812 592244
rect 442996 592080 443196 592244
rect 440650 591844 443196 592080
rect 440650 591680 442412 591844
rect 442596 591680 442812 591844
rect 442996 591680 443196 591844
rect 440650 591444 443196 591680
rect 440650 591280 442412 591444
rect 442596 591280 442812 591444
rect 442996 591280 443196 591444
rect 440650 591044 443196 591280
rect 440650 590880 442412 591044
rect 442596 590880 442822 591044
rect 443006 590880 443196 591044
rect 440650 590738 443196 590880
rect 446130 592148 448458 592380
rect 446130 591984 446212 592148
rect 446396 591984 446612 592148
rect 446796 591984 448458 592148
rect 446130 591748 448458 591984
rect 446130 591584 446212 591748
rect 446396 591584 446612 591748
rect 446796 591584 448458 591748
rect 446130 591348 448458 591584
rect 446130 591184 446212 591348
rect 446396 591184 446612 591348
rect 446796 591184 448458 591348
rect 446130 590948 448458 591184
rect 446130 590784 446212 590948
rect 446396 590784 446612 590948
rect 446796 590784 448458 590948
rect 446130 590716 448458 590784
rect 448998 592244 451596 592416
rect 448998 592080 450812 592244
rect 450996 592080 451212 592244
rect 451396 592080 451596 592244
rect 448998 591844 451596 592080
rect 448998 591680 450812 591844
rect 450996 591680 451212 591844
rect 451396 591680 451596 591844
rect 448998 591444 451596 591680
rect 448998 591280 450812 591444
rect 450996 591280 451212 591444
rect 451396 591280 451596 591444
rect 448998 591044 451596 591280
rect 448998 590880 450812 591044
rect 450996 590880 451222 591044
rect 451406 590880 451596 591044
rect 448998 590738 451596 590880
rect 448998 590736 449164 590738
rect 450322 590732 450740 590738
rect 438410 590704 440102 590716
rect 446810 590704 448458 590716
rect 440216 590212 440782 590254
rect 440216 590104 440260 590212
rect 440362 590104 440620 590212
rect 440722 590104 440782 590212
rect 440216 589972 440782 590104
rect 440216 589864 440260 589972
rect 440362 589864 440620 589972
rect 440722 589864 440782 589972
rect 440216 589824 440782 589864
rect 448544 590212 449110 590254
rect 448544 590104 448588 590212
rect 448690 590104 448948 590212
rect 449050 590104 449110 590212
rect 448544 589972 449110 590104
rect 448544 589864 448588 589972
rect 448690 589864 448948 589972
rect 449050 589864 449110 589972
rect 448544 589824 449110 589864
rect 406654 588654 408682 588724
rect 405388 588544 410080 588654
rect 405388 588304 405560 588544
rect 405868 588304 406160 588544
rect 406468 588304 406760 588544
rect 407068 588304 407360 588544
rect 407668 588304 407960 588544
rect 408268 588304 408560 588544
rect 408868 588304 409160 588544
rect 409468 588304 410080 588544
rect 405388 588224 410080 588304
rect 406654 587908 408682 588224
rect 404984 587696 405238 587706
rect 404984 587640 405006 587696
rect 405086 587640 405126 587696
rect 405206 587640 405238 587696
rect 404984 587596 405238 587640
rect 404984 587540 405006 587596
rect 405086 587540 405126 587596
rect 405206 587540 405238 587596
rect 404984 587510 405238 587540
rect 409968 587696 410212 587706
rect 409968 587640 409990 587696
rect 410070 587640 410110 587696
rect 410190 587640 410212 587696
rect 409968 587596 410212 587640
rect 409968 587540 409990 587596
rect 410070 587540 410110 587596
rect 410190 587540 410212 587596
rect 409968 587510 410212 587540
rect 404124 587104 404968 587106
rect 406648 587104 408678 587340
rect 404124 587030 410098 587104
rect 404124 586866 405398 587030
rect 405592 586866 405798 587030
rect 405992 586866 406198 587030
rect 406392 586866 406598 587030
rect 406792 586866 406998 587030
rect 407192 586866 407398 587030
rect 407592 586866 407798 587030
rect 407992 586866 408198 587030
rect 408392 586866 408598 587030
rect 408792 586866 408998 587030
rect 409192 586866 409398 587030
rect 409592 586866 409798 587030
rect 409992 586866 410098 587030
rect 404124 586790 410098 586866
rect 404124 586626 405398 586790
rect 405592 586626 405798 586790
rect 405992 586626 406198 586790
rect 406392 586626 406598 586790
rect 406792 586626 406998 586790
rect 407192 586626 407398 586790
rect 407592 586626 407798 586790
rect 407992 586626 408198 586790
rect 408392 586626 408598 586790
rect 408792 586626 408998 586790
rect 409192 586626 409398 586790
rect 409592 586626 409798 586790
rect 409992 586626 410098 586790
rect 404124 586572 410098 586626
rect 404124 586566 404968 586572
rect 404128 585078 404890 586566
rect 405230 586562 410092 586572
rect 405388 586344 410080 586454
rect 423906 586446 428284 586452
rect 438104 586450 440896 586452
rect 441242 586450 441936 586452
rect 433144 586446 441936 586450
rect 405388 586104 405560 586344
rect 405868 586104 406160 586344
rect 406468 586104 406760 586344
rect 407068 586104 407360 586344
rect 407668 586104 407960 586344
rect 408268 586104 408560 586344
rect 408868 586104 409160 586344
rect 409468 586104 410080 586344
rect 405388 586024 410080 586104
rect 416354 586336 417192 586444
rect 406642 585812 408672 586024
rect 416354 585948 416472 586336
rect 417092 586142 417192 586336
rect 423906 586394 441936 586446
rect 423906 586180 438974 586394
rect 441846 586214 441936 586394
rect 441846 586180 441958 586214
rect 417092 585948 418050 586142
rect 416354 585850 418050 585948
rect 417260 585844 418050 585850
rect 423906 586138 441958 586180
rect 423906 585792 424024 586138
rect 426680 586136 438282 586138
rect 426680 586132 433278 586136
rect 438896 586134 441958 586138
rect 426680 586126 428284 586132
rect 404984 585596 405258 585606
rect 404984 585540 405006 585596
rect 405086 585540 405126 585596
rect 405206 585540 405258 585596
rect 404984 585496 405258 585540
rect 404984 585440 405006 585496
rect 405086 585440 405126 585496
rect 405206 585440 405258 585496
rect 404984 585410 405258 585440
rect 409976 585596 410220 585606
rect 409976 585540 409998 585596
rect 410078 585540 410118 585596
rect 410198 585540 410220 585596
rect 409976 585496 410220 585540
rect 409976 585440 409998 585496
rect 410078 585440 410118 585496
rect 410198 585440 410220 585496
rect 409976 585410 410220 585440
rect 417068 585316 418090 585318
rect 404124 585076 405488 585078
rect 406642 585076 408668 585270
rect 416356 585216 418090 585316
rect 404124 585030 410092 585076
rect 404124 584866 405398 585030
rect 405592 584866 405798 585030
rect 405992 584866 406198 585030
rect 406392 584866 406598 585030
rect 406792 584866 406998 585030
rect 407192 584866 407398 585030
rect 407592 584866 407798 585030
rect 407992 584866 408198 585030
rect 408392 584866 408598 585030
rect 408792 584866 408998 585030
rect 409192 584866 409398 585030
rect 409592 584866 409798 585030
rect 409992 584866 410092 585030
rect 404124 584790 410092 584866
rect 404124 584626 405398 584790
rect 405592 584626 405798 584790
rect 405992 584626 406198 584790
rect 406392 584626 406598 584790
rect 406792 584626 406998 584790
rect 407192 584626 407398 584790
rect 407592 584626 407798 584790
rect 407992 584626 408198 584790
rect 408392 584626 408598 584790
rect 408792 584626 408998 584790
rect 409192 584626 409398 584790
rect 409592 584626 409798 584790
rect 409992 584626 410092 584790
rect 416356 584828 416474 585216
rect 417094 585020 418090 585216
rect 417094 584828 417188 585020
rect 417264 585018 418090 585020
rect 423906 585096 423996 585322
rect 426686 585096 450516 585098
rect 423906 585094 424068 585096
rect 424644 585094 450516 585096
rect 423906 585042 450516 585094
rect 416356 584730 417188 584828
rect 423906 584840 447368 585042
rect 450242 584840 450516 585042
rect 423906 584792 450516 584840
rect 426686 584790 450516 584792
rect 404124 584538 410092 584626
rect 404128 584534 404890 584538
rect 405236 582858 410092 584538
rect 405234 581174 410096 582858
rect 405234 580628 405622 581174
rect 406400 580628 406822 581174
rect 407600 580628 408022 581174
rect 408800 580628 409222 581174
rect 410000 580628 410096 581174
rect 405234 580228 410096 580628
<< via1 >>
rect 119008 695372 119292 695430
rect 119008 695204 119058 695372
rect 119058 695204 119246 695372
rect 119246 695204 119292 695372
rect 119008 695156 119292 695204
rect 120660 694918 121252 695446
rect 121760 694918 122352 695446
rect 122860 694918 123452 695446
rect 123960 694918 124552 695446
rect 126230 695110 126562 695464
rect 415392 691208 415494 691316
rect 415752 691208 415854 691316
rect 415392 690968 415494 691076
rect 415752 690968 415854 691076
rect 467296 691308 467398 691416
rect 467656 691308 467758 691416
rect 467296 691068 467398 691176
rect 467656 691068 467758 691176
rect 569260 691308 569362 691416
rect 569620 691308 569722 691416
rect 569260 691068 569362 691176
rect 569620 691068 569722 691176
rect 571002 689284 571242 689592
rect 413812 688212 413996 688376
rect 414212 688212 414396 688376
rect 413812 687812 413996 687976
rect 414212 687812 414396 687976
rect 67008 687402 67292 687430
rect 67008 687178 67028 687402
rect 67028 687178 67270 687402
rect 67270 687178 67292 687402
rect 67008 687156 67292 687178
rect 68660 686918 69252 687446
rect 69760 686918 70352 687446
rect 70860 686918 71452 687446
rect 71960 686918 72552 687446
rect 74230 687110 74562 687464
rect 413812 687412 413996 687576
rect 414212 687412 414396 687576
rect 413812 687012 413996 687176
rect 414212 687012 414396 687176
rect 416278 688212 416396 688376
rect 416612 688212 416796 688376
rect 416278 687812 416396 687976
rect 416612 687812 416796 687976
rect 416278 687412 416396 687576
rect 416612 687412 416796 687576
rect 416278 687012 416396 687176
rect 416622 687012 416806 687176
rect 465812 688212 465996 688376
rect 466212 688212 466396 688376
rect 465812 687812 465996 687976
rect 466212 687812 466396 687976
rect 465812 687412 465996 687576
rect 466212 687412 466396 687576
rect 465812 687012 465996 687176
rect 466212 687012 466396 687176
rect 571002 688684 571242 688992
rect 468212 688212 468396 688376
rect 468612 688212 468796 688376
rect 468212 687812 468396 687976
rect 468612 687812 468796 687976
rect 468212 687412 468396 687576
rect 468612 687412 468796 687576
rect 468212 687012 468396 687176
rect 468622 687012 468806 687176
rect 568212 688212 568396 688376
rect 568612 688212 568796 688376
rect 568212 687812 568396 687976
rect 568612 687812 568796 687976
rect 568212 687412 568396 687576
rect 568612 687412 568796 687576
rect 568212 687012 568396 687176
rect 568622 687012 568806 687176
rect 571002 688084 571242 688392
rect 571002 687484 571242 687792
rect 571002 686884 571242 687192
rect 571002 686284 571242 686592
rect 571002 685684 571242 685992
rect 415606 685408 415708 685516
rect 415966 685408 416068 685516
rect 415606 685168 415708 685276
rect 415966 685168 416068 685276
rect 467190 685404 467292 685512
rect 467550 685404 467652 685512
rect 467190 685164 467292 685272
rect 467550 685164 467652 685272
rect 569260 683708 569362 683816
rect 569620 683708 569722 683816
rect 569260 683468 569362 683576
rect 569620 683468 569722 683576
rect 70580 674824 70682 674932
rect 70940 674824 71042 674932
rect 70580 674584 70682 674692
rect 70940 674584 71042 674692
rect 122568 674866 122670 674974
rect 122928 674866 123030 674974
rect 122568 674626 122670 674734
rect 122928 674626 123030 674734
rect 70008 673458 70292 673732
rect 71368 673402 71700 673756
rect 121808 673220 122092 673494
rect 123302 673110 123634 673464
rect 70570 672224 70672 672332
rect 70930 672224 71032 672332
rect 70570 671984 70672 672092
rect 70930 671984 71032 672092
rect 122558 672266 122660 672374
rect 122918 672266 123020 672374
rect 122558 672026 122660 672134
rect 122918 672026 123020 672134
rect 440252 593576 440354 593684
rect 440612 593576 440714 593684
rect 440252 593336 440354 593444
rect 440612 593336 440714 593444
rect 448600 593608 448702 593716
rect 448960 593608 449062 593716
rect 448600 593368 448702 593476
rect 448960 593368 449062 593476
rect 437812 591984 437996 592148
rect 438212 591984 438396 592148
rect 437812 591584 437996 591748
rect 438212 591584 438396 591748
rect 437812 591184 437996 591348
rect 438212 591184 438396 591348
rect 437812 590784 437996 590948
rect 438212 590784 438396 590948
rect 442412 592080 442596 592244
rect 442812 592080 442996 592244
rect 442412 591680 442596 591844
rect 442812 591680 442996 591844
rect 442412 591280 442596 591444
rect 442812 591280 442996 591444
rect 442412 590880 442596 591044
rect 442822 590880 443006 591044
rect 446212 591984 446396 592148
rect 446612 591984 446796 592148
rect 446212 591584 446396 591748
rect 446612 591584 446796 591748
rect 446212 591184 446396 591348
rect 446612 591184 446796 591348
rect 446212 590784 446396 590948
rect 446612 590784 446796 590948
rect 450812 592080 450996 592244
rect 451212 592080 451396 592244
rect 450812 591680 450996 591844
rect 451212 591680 451396 591844
rect 450812 591280 450996 591444
rect 451212 591280 451396 591444
rect 450812 590880 450996 591044
rect 451222 590880 451406 591044
rect 440260 590104 440362 590212
rect 440620 590104 440722 590212
rect 440260 589864 440362 589972
rect 440620 589864 440722 589972
rect 448588 590104 448690 590212
rect 448948 590104 449050 590212
rect 448588 589864 448690 589972
rect 448948 589864 449050 589972
rect 405560 588304 405868 588544
rect 406160 588304 406468 588544
rect 406760 588304 407068 588544
rect 407360 588304 407668 588544
rect 407960 588304 408268 588544
rect 408560 588304 408868 588544
rect 409160 588304 409468 588544
rect 405006 587640 405086 587696
rect 405126 587640 405206 587696
rect 405006 587540 405086 587596
rect 405126 587540 405206 587596
rect 409990 587640 410070 587696
rect 410110 587640 410190 587696
rect 409990 587540 410070 587596
rect 410110 587540 410190 587596
rect 405560 586104 405868 586344
rect 406160 586104 406468 586344
rect 406760 586104 407068 586344
rect 407360 586104 407668 586344
rect 407960 586104 408268 586344
rect 408560 586104 408868 586344
rect 409160 586104 409468 586344
rect 416472 585948 417092 586336
rect 438974 586180 441846 586394
rect 405006 585540 405086 585596
rect 405126 585540 405206 585596
rect 405006 585440 405086 585496
rect 405126 585440 405206 585496
rect 409998 585540 410078 585596
rect 410118 585540 410198 585596
rect 409998 585440 410078 585496
rect 410118 585440 410198 585496
rect 416474 584828 417094 585216
rect 447368 584840 450242 585042
rect 405622 580628 406400 581174
rect 406822 580628 407600 581174
rect 408022 580628 408800 581174
rect 409222 580628 410000 581174
<< metal2 >>
rect 118982 695430 119314 695454
rect 118982 695156 119008 695430
rect 119292 695156 119314 695430
rect 118982 695134 119314 695156
rect 120228 695446 124764 696194
rect 120228 694918 120660 695446
rect 121252 694918 121760 695446
rect 122352 694918 122860 695446
rect 123452 694918 123960 695446
rect 124552 694918 124764 695446
rect 126152 695464 126622 695524
rect 126152 695110 126230 695464
rect 126562 695110 126622 695464
rect 126152 695052 126622 695110
rect 120228 694328 124764 694918
rect 467252 691416 467818 691454
rect 415348 691316 415914 691358
rect 415348 691208 415392 691316
rect 415494 691208 415752 691316
rect 415854 691208 415914 691316
rect 415348 691076 415914 691208
rect 415348 690968 415392 691076
rect 415494 690968 415752 691076
rect 415854 690968 415914 691076
rect 467252 691308 467296 691416
rect 467398 691308 467656 691416
rect 467758 691308 467818 691416
rect 467252 691176 467818 691308
rect 467252 691068 467296 691176
rect 467398 691068 467656 691176
rect 467758 691068 467818 691176
rect 467252 691026 467818 691068
rect 569216 691416 569782 691454
rect 569216 691308 569260 691416
rect 569362 691308 569620 691416
rect 569722 691308 569782 691416
rect 569216 691176 569782 691308
rect 569216 691068 569260 691176
rect 569362 691068 569620 691176
rect 569722 691068 569782 691176
rect 569216 691028 569782 691068
rect 415348 690926 415914 690968
rect 570922 689592 571352 689764
rect 570922 689284 571002 689592
rect 571242 689284 571352 689592
rect 570922 688992 571352 689284
rect 570922 688684 571002 688992
rect 571242 688684 571352 688992
rect 413730 688376 414462 688608
rect 413730 688212 413812 688376
rect 413996 688212 414212 688376
rect 414396 688212 414462 688376
rect 66982 687430 67314 687454
rect 66982 687156 67008 687430
rect 67292 687156 67314 687430
rect 66982 687134 67314 687156
rect 68228 687446 72764 688194
rect 413730 687976 414462 688212
rect 413730 687812 413812 687976
rect 413996 687812 414212 687976
rect 414396 687812 414462 687976
rect 413730 687576 414462 687812
rect 68228 686918 68660 687446
rect 69252 686918 69760 687446
rect 70352 686918 70860 687446
rect 71452 686918 71960 687446
rect 72552 686918 72764 687446
rect 74152 687464 74622 687524
rect 74152 687110 74230 687464
rect 74562 687110 74622 687464
rect 74152 687052 74622 687110
rect 413730 687412 413812 687576
rect 413996 687412 414212 687576
rect 414396 687412 414462 687576
rect 413730 687176 414462 687412
rect 413730 687012 413812 687176
rect 413996 687012 414212 687176
rect 414396 687012 414462 687176
rect 413730 686944 414462 687012
rect 416130 688376 416866 688598
rect 416130 688212 416212 688376
rect 416396 688212 416612 688376
rect 416796 688212 416866 688376
rect 416130 687976 416866 688212
rect 416130 687812 416212 687976
rect 416396 687812 416612 687976
rect 416796 687812 416866 687976
rect 416130 687576 416866 687812
rect 416130 687412 416212 687576
rect 416396 687412 416612 687576
rect 416796 687412 416866 687576
rect 416130 687176 416866 687412
rect 416130 687012 416212 687176
rect 416396 687012 416622 687176
rect 416806 687012 416866 687176
rect 416130 686944 416866 687012
rect 465730 688376 466466 688608
rect 465730 688212 465812 688376
rect 465996 688212 466212 688376
rect 466396 688212 466466 688376
rect 465730 687976 466466 688212
rect 465730 687812 465812 687976
rect 465996 687812 466212 687976
rect 466396 687812 466466 687976
rect 465730 687576 466466 687812
rect 465730 687412 465812 687576
rect 465996 687412 466212 687576
rect 466396 687412 466466 687576
rect 465730 687176 466466 687412
rect 465730 687012 465812 687176
rect 465996 687012 466212 687176
rect 466396 687012 466466 687176
rect 465730 686944 466466 687012
rect 468130 688376 468866 688598
rect 468130 688212 468212 688376
rect 468396 688212 468612 688376
rect 468796 688212 468866 688376
rect 468130 687976 468866 688212
rect 468130 687812 468212 687976
rect 468396 687812 468612 687976
rect 468796 687812 468866 687976
rect 468130 687576 468866 687812
rect 468130 687412 468212 687576
rect 468396 687412 468612 687576
rect 468796 687412 468866 687576
rect 468130 687176 468866 687412
rect 468130 687012 468212 687176
rect 468396 687012 468622 687176
rect 468806 687012 468866 687176
rect 468130 686944 468866 687012
rect 568130 688376 568866 688598
rect 568130 688212 568212 688376
rect 568396 688212 568612 688376
rect 568796 688212 568866 688376
rect 568130 687976 568866 688212
rect 568130 687812 568212 687976
rect 568396 687812 568612 687976
rect 568796 687812 568866 687976
rect 568130 687576 568866 687812
rect 568130 687412 568212 687576
rect 568396 687412 568612 687576
rect 568796 687412 568866 687576
rect 568130 687176 568866 687412
rect 568130 687012 568212 687176
rect 568396 687012 568622 687176
rect 568806 687012 568866 687176
rect 568130 686944 568866 687012
rect 570922 688392 571352 688684
rect 570922 688084 571002 688392
rect 571242 688084 571352 688392
rect 570922 687792 571352 688084
rect 570922 687484 571002 687792
rect 571242 687484 571352 687792
rect 570922 687192 571352 687484
rect 68228 686328 72764 686918
rect 570922 686884 571002 687192
rect 571242 686884 571352 687192
rect 570922 686592 571352 686884
rect 570922 686284 571002 686592
rect 571242 686284 571352 686592
rect 570922 685992 571352 686284
rect 570922 685684 571002 685992
rect 571242 685684 571352 685992
rect 415562 685516 416128 685558
rect 415562 685408 415606 685516
rect 415708 685408 415966 685516
rect 416068 685408 416128 685516
rect 415562 685276 416128 685408
rect 415562 685168 415606 685276
rect 415708 685168 415966 685276
rect 416068 685168 416128 685276
rect 415562 685126 416128 685168
rect 467146 685554 467272 685580
rect 467146 685512 467712 685554
rect 467146 685404 467190 685512
rect 467292 685404 467550 685512
rect 467652 685404 467712 685512
rect 467146 685272 467712 685404
rect 467146 685164 467190 685272
rect 467292 685164 467550 685272
rect 467652 685164 467712 685272
rect 467146 685122 467712 685164
rect 570922 685072 571352 685684
rect 569216 683816 569782 683852
rect 569216 683814 569260 683816
rect 569362 683814 569620 683816
rect 569216 683466 569256 683814
rect 569722 683466 569782 683816
rect 569216 683434 569782 683466
rect 122524 674974 123090 675016
rect 70536 674932 71102 674974
rect 70536 674824 70580 674932
rect 70682 674824 70940 674932
rect 71042 674824 71102 674932
rect 70536 674692 71102 674824
rect 70536 674584 70580 674692
rect 70682 674584 70940 674692
rect 71042 674584 71102 674692
rect 122524 674866 122568 674974
rect 122670 674866 122928 674974
rect 123030 674866 123090 674974
rect 122524 674734 123090 674866
rect 122524 674626 122568 674734
rect 122670 674626 122928 674734
rect 123030 674626 123090 674734
rect 122524 674586 123090 674626
rect 70536 674544 71102 674584
rect 71290 673756 71760 673816
rect 69982 673732 70314 673756
rect 69982 673458 70008 673732
rect 70292 673458 70314 673732
rect 69982 673436 70314 673458
rect 71290 673402 71368 673756
rect 71700 673402 71760 673756
rect 71290 673344 71760 673402
rect 121782 673494 122114 673518
rect 121782 673220 121808 673494
rect 122092 673220 122114 673494
rect 121782 673198 122114 673220
rect 123224 673464 123694 673524
rect 123224 673110 123302 673464
rect 123634 673110 123694 673464
rect 123224 673052 123694 673110
rect 122514 672374 123080 672416
rect 70526 672332 71092 672374
rect 70526 672224 70570 672332
rect 70672 672224 70930 672332
rect 71032 672224 71092 672332
rect 70526 672092 71092 672224
rect 70526 671984 70570 672092
rect 70672 671984 70930 672092
rect 71032 671984 71092 672092
rect 122514 672266 122558 672374
rect 122660 672266 122918 672374
rect 123020 672266 123080 672374
rect 122514 672134 123080 672266
rect 122514 672026 122558 672134
rect 122660 672026 122918 672134
rect 123020 672026 123080 672134
rect 122514 671986 123080 672026
rect 70526 671944 71092 671984
rect 440208 593684 440774 593726
rect 440208 593576 440252 593684
rect 440354 593576 440612 593684
rect 440714 593576 440774 593684
rect 440208 593444 440774 593576
rect 440208 593336 440252 593444
rect 440354 593336 440612 593444
rect 440714 593336 440774 593444
rect 440208 593296 440774 593336
rect 448556 593716 449122 593758
rect 448556 593608 448600 593716
rect 448702 593608 448960 593716
rect 449062 593608 449122 593716
rect 448556 593476 449122 593608
rect 448556 593368 448600 593476
rect 448702 593368 448960 593476
rect 449062 593368 449122 593476
rect 448556 593328 449122 593368
rect 437730 592148 438466 592380
rect 437730 591984 437812 592148
rect 437996 591984 438212 592148
rect 438396 591984 438466 592148
rect 437730 591748 438466 591984
rect 437730 591584 437812 591748
rect 437996 591584 438212 591748
rect 438396 591584 438466 591748
rect 437730 591348 438466 591584
rect 437730 591184 437812 591348
rect 437996 591184 438212 591348
rect 438396 591184 438466 591348
rect 437730 590948 438466 591184
rect 437730 590784 437812 590948
rect 437996 590784 438212 590948
rect 438396 590784 438466 590948
rect 442330 592244 443066 592420
rect 442330 592080 442412 592244
rect 442596 592080 442812 592244
rect 442996 592080 443066 592244
rect 442330 591844 443066 592080
rect 442330 591680 442412 591844
rect 442596 591680 442812 591844
rect 442996 591680 443066 591844
rect 442330 591444 443066 591680
rect 442330 591280 442412 591444
rect 442596 591280 442812 591444
rect 442996 591280 443066 591444
rect 442330 591044 443066 591280
rect 442330 590880 442412 591044
rect 442596 590880 442822 591044
rect 443006 590880 443066 591044
rect 442330 590812 443066 590880
rect 446130 592148 446866 592380
rect 446130 591984 446212 592148
rect 446396 591984 446612 592148
rect 446796 591984 446866 592148
rect 446130 591748 446866 591984
rect 446130 591584 446212 591748
rect 446396 591584 446612 591748
rect 446796 591584 446866 591748
rect 446130 591348 446866 591584
rect 446130 591184 446212 591348
rect 446396 591184 446612 591348
rect 446796 591184 446866 591348
rect 446130 590948 446866 591184
rect 437730 590716 438466 590784
rect 446130 590784 446212 590948
rect 446396 590784 446612 590948
rect 446796 590784 446866 590948
rect 450730 592244 451466 592420
rect 450730 592080 450812 592244
rect 450996 592080 451212 592244
rect 451396 592080 451466 592244
rect 450730 591844 451466 592080
rect 450730 591680 450812 591844
rect 450996 591680 451212 591844
rect 451396 591680 451466 591844
rect 450730 591444 451466 591680
rect 450730 591280 450812 591444
rect 450996 591280 451212 591444
rect 451396 591280 451466 591444
rect 450730 591044 451466 591280
rect 450730 590880 450812 591044
rect 450996 590880 451222 591044
rect 451406 590880 451466 591044
rect 450730 590812 451466 590880
rect 446130 590716 446866 590784
rect 440216 590212 440782 590254
rect 440216 590104 440260 590212
rect 440362 590104 440620 590212
rect 440722 590104 440782 590212
rect 440216 589972 440782 590104
rect 440216 589864 440260 589972
rect 440362 589864 440620 589972
rect 440722 589864 440782 589972
rect 440216 589824 440782 589864
rect 448544 590212 449110 590254
rect 448544 590104 448588 590212
rect 448690 590104 448948 590212
rect 449050 590104 449110 590212
rect 448544 589972 449110 590104
rect 448544 589864 448588 589972
rect 448690 589864 448948 589972
rect 449050 589864 449110 589972
rect 448544 589824 449110 589864
rect 405388 588544 410080 588654
rect 405388 588304 405560 588544
rect 405868 588304 406160 588544
rect 406468 588304 406760 588544
rect 407068 588304 407360 588544
rect 407668 588304 407960 588544
rect 408268 588304 408560 588544
rect 408868 588304 409160 588544
rect 409468 588304 410080 588544
rect 405388 588224 410080 588304
rect 404984 587696 405238 587706
rect 404984 587640 405006 587696
rect 405086 587640 405126 587696
rect 405206 587640 405238 587696
rect 404984 587596 405238 587640
rect 404984 587540 405006 587596
rect 405086 587540 405126 587596
rect 405206 587540 405238 587596
rect 404984 587510 405238 587540
rect 409968 587696 410212 587706
rect 409968 587640 409990 587696
rect 410070 587640 410110 587696
rect 410190 587640 410212 587696
rect 409968 587596 410212 587640
rect 409968 587540 409990 587596
rect 410070 587540 410110 587596
rect 410190 587540 410212 587596
rect 409968 587510 410212 587540
rect 405388 586344 410080 586454
rect 405388 586104 405560 586344
rect 405868 586104 406160 586344
rect 406468 586104 406760 586344
rect 407068 586104 407360 586344
rect 407668 586104 407960 586344
rect 408268 586104 408560 586344
rect 408868 586104 409160 586344
rect 409468 586104 410080 586344
rect 405388 586024 410080 586104
rect 416354 586336 417192 586444
rect 416354 585948 416472 586336
rect 417092 585948 417192 586336
rect 438926 586394 441902 586434
rect 438926 586180 438974 586394
rect 441846 586180 441902 586394
rect 438926 586136 441902 586180
rect 416354 585850 417192 585948
rect 404984 585596 405258 585606
rect 404984 585540 405006 585596
rect 405086 585540 405126 585596
rect 405206 585540 405258 585596
rect 404984 585496 405258 585540
rect 404984 585440 405006 585496
rect 405086 585440 405126 585496
rect 405206 585440 405258 585496
rect 404984 585410 405258 585440
rect 409976 585596 410220 585606
rect 409976 585540 409998 585596
rect 410078 585540 410118 585596
rect 410198 585540 410220 585596
rect 409976 585496 410220 585540
rect 409976 585440 409998 585496
rect 410078 585440 410118 585496
rect 410198 585440 410220 585496
rect 409976 585410 410220 585440
rect 416356 585216 417188 585316
rect 416356 584828 416474 585216
rect 417094 584828 417188 585216
rect 416356 584730 417188 584828
rect 447352 585042 450258 585064
rect 447352 584840 447368 585042
rect 450242 584840 450258 585042
rect 447352 584820 450258 584840
rect 405234 581174 410146 581588
rect 405234 580628 405622 581174
rect 406400 580628 406822 581174
rect 407600 580628 408022 581174
rect 408800 580628 409222 581174
rect 410000 580628 410146 581174
rect 405234 580232 410146 580628
rect 524 -800 636 480
rect 1706 -800 1818 480
rect 2888 -800 3000 480
rect 4070 -800 4182 480
rect 5252 -800 5364 480
rect 6434 -800 6546 480
rect 7616 -800 7728 480
rect 8798 -800 8910 480
rect 9980 -800 10092 480
rect 11162 -800 11274 480
rect 12344 -800 12456 480
rect 13526 -800 13638 480
rect 14708 -800 14820 480
rect 15890 -800 16002 480
rect 17072 -800 17184 480
rect 18254 -800 18366 480
rect 19436 -800 19548 480
rect 20618 -800 20730 480
rect 21800 -800 21912 480
rect 22982 -800 23094 480
rect 24164 -800 24276 480
rect 25346 -800 25458 480
rect 26528 -800 26640 480
rect 27710 -800 27822 480
rect 28892 -800 29004 480
rect 30074 -800 30186 480
rect 31256 -800 31368 480
rect 32438 -800 32550 480
rect 33620 -800 33732 480
rect 34802 -800 34914 480
rect 35984 -800 36096 480
rect 37166 -800 37278 480
rect 38348 -800 38460 480
rect 39530 -800 39642 480
rect 40712 -800 40824 480
rect 41894 -800 42006 480
rect 43076 -800 43188 480
rect 44258 -800 44370 480
rect 45440 -800 45552 480
rect 46622 -800 46734 480
rect 47804 -800 47916 480
rect 48986 -800 49098 480
rect 50168 -800 50280 480
rect 51350 -800 51462 480
rect 52532 -800 52644 480
rect 53714 -800 53826 480
rect 54896 -800 55008 480
rect 56078 -800 56190 480
rect 57260 -800 57372 480
rect 58442 -800 58554 480
rect 59624 -800 59736 480
rect 60806 -800 60918 480
rect 61988 -800 62100 480
rect 63170 -800 63282 480
rect 64352 -800 64464 480
rect 65534 -800 65646 480
rect 66716 -800 66828 480
rect 67898 -800 68010 480
rect 69080 -800 69192 480
rect 70262 -800 70374 480
rect 71444 -800 71556 480
rect 72626 -800 72738 480
rect 73808 -800 73920 480
rect 74990 -800 75102 480
rect 76172 -800 76284 480
rect 77354 -800 77466 480
rect 78536 -800 78648 480
rect 79718 -800 79830 480
rect 80900 -800 81012 480
rect 82082 -800 82194 480
rect 83264 -800 83376 480
rect 84446 -800 84558 480
rect 85628 -800 85740 480
rect 86810 -800 86922 480
rect 87992 -800 88104 480
rect 89174 -800 89286 480
rect 90356 -800 90468 480
rect 91538 -800 91650 480
rect 92720 -800 92832 480
rect 93902 -800 94014 480
rect 95084 -800 95196 480
rect 96266 -800 96378 480
rect 97448 -800 97560 480
rect 98630 -800 98742 480
rect 99812 -800 99924 480
rect 100994 -800 101106 480
rect 102176 -800 102288 480
rect 103358 -800 103470 480
rect 104540 -800 104652 480
rect 105722 -800 105834 480
rect 106904 -800 107016 480
rect 108086 -800 108198 480
rect 109268 -800 109380 480
rect 110450 -800 110562 480
rect 111632 -800 111744 480
rect 112814 -800 112926 480
rect 113996 -800 114108 480
rect 115178 -800 115290 480
rect 116360 -800 116472 480
rect 117542 -800 117654 480
rect 118724 -800 118836 480
rect 119906 -800 120018 480
rect 121088 -800 121200 480
rect 122270 -800 122382 480
rect 123452 -800 123564 480
rect 124634 -800 124746 480
rect 125816 -800 125928 480
rect 126998 -800 127110 480
rect 128180 -800 128292 480
rect 129362 -800 129474 480
rect 130544 -800 130656 480
rect 131726 -800 131838 480
rect 132908 -800 133020 480
rect 134090 -800 134202 480
rect 135272 -800 135384 480
rect 136454 -800 136566 480
rect 137636 -800 137748 480
rect 138818 -800 138930 480
rect 140000 -800 140112 480
rect 141182 -800 141294 480
rect 142364 -800 142476 480
rect 143546 -800 143658 480
rect 144728 -800 144840 480
rect 145910 -800 146022 480
rect 147092 -800 147204 480
rect 148274 -800 148386 480
rect 149456 -800 149568 480
rect 150638 -800 150750 480
rect 151820 -800 151932 480
rect 153002 -800 153114 480
rect 154184 -800 154296 480
rect 155366 -800 155478 480
rect 156548 -800 156660 480
rect 157730 -800 157842 480
rect 158912 -800 159024 480
rect 160094 -800 160206 480
rect 161276 -800 161388 480
rect 162458 -800 162570 480
rect 163640 -800 163752 480
rect 164822 -800 164934 480
rect 166004 -800 166116 480
rect 167186 -800 167298 480
rect 168368 -800 168480 480
rect 169550 -800 169662 480
rect 170732 -800 170844 480
rect 171914 -800 172026 480
rect 173096 -800 173208 480
rect 174278 -800 174390 480
rect 175460 -800 175572 480
rect 176642 -800 176754 480
rect 177824 -800 177936 480
rect 179006 -800 179118 480
rect 180188 -800 180300 480
rect 181370 -800 181482 480
rect 182552 -800 182664 480
rect 183734 -800 183846 480
rect 184916 -800 185028 480
rect 186098 -800 186210 480
rect 187280 -800 187392 480
rect 188462 -800 188574 480
rect 189644 -800 189756 480
rect 190826 -800 190938 480
rect 192008 -800 192120 480
rect 193190 -800 193302 480
rect 194372 -800 194484 480
rect 195554 -800 195666 480
rect 196736 -800 196848 480
rect 197918 -800 198030 480
rect 199100 -800 199212 480
rect 200282 -800 200394 480
rect 201464 -800 201576 480
rect 202646 -800 202758 480
rect 203828 -800 203940 480
rect 205010 -800 205122 480
rect 206192 -800 206304 480
rect 207374 -800 207486 480
rect 208556 -800 208668 480
rect 209738 -800 209850 480
rect 210920 -800 211032 480
rect 212102 -800 212214 480
rect 213284 -800 213396 480
rect 214466 -800 214578 480
rect 215648 -800 215760 480
rect 216830 -800 216942 480
rect 218012 -800 218124 480
rect 219194 -800 219306 480
rect 220376 -800 220488 480
rect 221558 -800 221670 480
rect 222740 -800 222852 480
rect 223922 -800 224034 480
rect 225104 -800 225216 480
rect 226286 -800 226398 480
rect 227468 -800 227580 480
rect 228650 -800 228762 480
rect 229832 -800 229944 480
rect 231014 -800 231126 480
rect 232196 -800 232308 480
rect 233378 -800 233490 480
rect 234560 -800 234672 480
rect 235742 -800 235854 480
rect 236924 -800 237036 480
rect 238106 -800 238218 480
rect 239288 -800 239400 480
rect 240470 -800 240582 480
rect 241652 -800 241764 480
rect 242834 -800 242946 480
rect 244016 -800 244128 480
rect 245198 -800 245310 480
rect 246380 -800 246492 480
rect 247562 -800 247674 480
rect 248744 -800 248856 480
rect 249926 -800 250038 480
rect 251108 -800 251220 480
rect 252290 -800 252402 480
rect 253472 -800 253584 480
rect 254654 -800 254766 480
rect 255836 -800 255948 480
rect 257018 -800 257130 480
rect 258200 -800 258312 480
rect 259382 -800 259494 480
rect 260564 -800 260676 480
rect 261746 -800 261858 480
rect 262928 -800 263040 480
rect 264110 -800 264222 480
rect 265292 -800 265404 480
rect 266474 -800 266586 480
rect 267656 -800 267768 480
rect 268838 -800 268950 480
rect 270020 -800 270132 480
rect 271202 -800 271314 480
rect 272384 -800 272496 480
rect 273566 -800 273678 480
rect 274748 -800 274860 480
rect 275930 -800 276042 480
rect 277112 -800 277224 480
rect 278294 -800 278406 480
rect 279476 -800 279588 480
rect 280658 -800 280770 480
rect 281840 -800 281952 480
rect 283022 -800 283134 480
rect 284204 -800 284316 480
rect 285386 -800 285498 480
rect 286568 -800 286680 480
rect 287750 -800 287862 480
rect 288932 -800 289044 480
rect 290114 -800 290226 480
rect 291296 -800 291408 480
rect 292478 -800 292590 480
rect 293660 -800 293772 480
rect 294842 -800 294954 480
rect 296024 -800 296136 480
rect 297206 -800 297318 480
rect 298388 -800 298500 480
rect 299570 -800 299682 480
rect 300752 -800 300864 480
rect 301934 -800 302046 480
rect 303116 -800 303228 480
rect 304298 -800 304410 480
rect 305480 -800 305592 480
rect 306662 -800 306774 480
rect 307844 -800 307956 480
rect 309026 -800 309138 480
rect 310208 -800 310320 480
rect 311390 -800 311502 480
rect 312572 -800 312684 480
rect 313754 -800 313866 480
rect 314936 -800 315048 480
rect 316118 -800 316230 480
rect 317300 -800 317412 480
rect 318482 -800 318594 480
rect 319664 -800 319776 480
rect 320846 -800 320958 480
rect 322028 -800 322140 480
rect 323210 -800 323322 480
rect 324392 -800 324504 480
rect 325574 -800 325686 480
rect 326756 -800 326868 480
rect 327938 -800 328050 480
rect 329120 -800 329232 480
rect 330302 -800 330414 480
rect 331484 -800 331596 480
rect 332666 -800 332778 480
rect 333848 -800 333960 480
rect 335030 -800 335142 480
rect 336212 -800 336324 480
rect 337394 -800 337506 480
rect 338576 -800 338688 480
rect 339758 -800 339870 480
rect 340940 -800 341052 480
rect 342122 -800 342234 480
rect 343304 -800 343416 480
rect 344486 -800 344598 480
rect 345668 -800 345780 480
rect 346850 -800 346962 480
rect 348032 -800 348144 480
rect 349214 -800 349326 480
rect 350396 -800 350508 480
rect 351578 -800 351690 480
rect 352760 -800 352872 480
rect 353942 -800 354054 480
rect 355124 -800 355236 480
rect 356306 -800 356418 480
rect 357488 -800 357600 480
rect 358670 -800 358782 480
rect 359852 -800 359964 480
rect 361034 -800 361146 480
rect 362216 -800 362328 480
rect 363398 -800 363510 480
rect 364580 -800 364692 480
rect 365762 -800 365874 480
rect 366944 -800 367056 480
rect 368126 -800 368238 480
rect 369308 -800 369420 480
rect 370490 -800 370602 480
rect 371672 -800 371784 480
rect 372854 -800 372966 480
rect 374036 -800 374148 480
rect 375218 -800 375330 480
rect 376400 -800 376512 480
rect 377582 -800 377694 480
rect 378764 -800 378876 480
rect 379946 -800 380058 480
rect 381128 -800 381240 480
rect 382310 -800 382422 480
rect 383492 -800 383604 480
rect 384674 -800 384786 480
rect 385856 -800 385968 480
rect 387038 -800 387150 480
rect 388220 -800 388332 480
rect 389402 -800 389514 480
rect 390584 -800 390696 480
rect 391766 -800 391878 480
rect 392948 -800 393060 480
rect 394130 -800 394242 480
rect 395312 -800 395424 480
rect 396494 -800 396606 480
rect 397676 -800 397788 480
rect 398858 -800 398970 480
rect 400040 -800 400152 480
rect 401222 -800 401334 480
rect 402404 -800 402516 480
rect 403586 -800 403698 480
rect 404768 -800 404880 480
rect 405950 -800 406062 480
rect 407132 -800 407244 480
rect 408314 -800 408426 480
rect 409496 -800 409608 480
rect 410678 -800 410790 480
rect 411860 -800 411972 480
rect 413042 -800 413154 480
rect 414224 -800 414336 480
rect 415406 -800 415518 480
rect 416588 -800 416700 480
rect 417770 -800 417882 480
rect 418952 -800 419064 480
rect 420134 -800 420246 480
rect 421316 -800 421428 480
rect 422498 -800 422610 480
rect 423680 -800 423792 480
rect 424862 -800 424974 480
rect 426044 -800 426156 480
rect 427226 -800 427338 480
rect 428408 -800 428520 480
rect 429590 -800 429702 480
rect 430772 -800 430884 480
rect 431954 -800 432066 480
rect 433136 -800 433248 480
rect 434318 -800 434430 480
rect 435500 -800 435612 480
rect 436682 -800 436794 480
rect 437864 -800 437976 480
rect 439046 -800 439158 480
rect 440228 -800 440340 480
rect 441410 -800 441522 480
rect 442592 -800 442704 480
rect 443774 -800 443886 480
rect 444956 -800 445068 480
rect 446138 -800 446250 480
rect 447320 -800 447432 480
rect 448502 -800 448614 480
rect 449684 -800 449796 480
rect 450866 -800 450978 480
rect 452048 -800 452160 480
rect 453230 -800 453342 480
rect 454412 -800 454524 480
rect 455594 -800 455706 480
rect 456776 -800 456888 480
rect 457958 -800 458070 480
rect 459140 -800 459252 480
rect 460322 -800 460434 480
rect 461504 -800 461616 480
rect 462686 -800 462798 480
rect 463868 -800 463980 480
rect 465050 -800 465162 480
rect 466232 -800 466344 480
rect 467414 -800 467526 480
rect 468596 -800 468708 480
rect 469778 -800 469890 480
rect 470960 -800 471072 480
rect 472142 -800 472254 480
rect 473324 -800 473436 480
rect 474506 -800 474618 480
rect 475688 -800 475800 480
rect 476870 -800 476982 480
rect 478052 -800 478164 480
rect 479234 -800 479346 480
rect 480416 -800 480528 480
rect 481598 -800 481710 480
rect 482780 -800 482892 480
rect 483962 -800 484074 480
rect 485144 -800 485256 480
rect 486326 -800 486438 480
rect 487508 -800 487620 480
rect 488690 -800 488802 480
rect 489872 -800 489984 480
rect 491054 -800 491166 480
rect 492236 -800 492348 480
rect 493418 -800 493530 480
rect 494600 -800 494712 480
rect 495782 -800 495894 480
rect 496964 -800 497076 480
rect 498146 -800 498258 480
rect 499328 -800 499440 480
rect 500510 -800 500622 480
rect 501692 -800 501804 480
rect 502874 -800 502986 480
rect 504056 -800 504168 480
rect 505238 -800 505350 480
rect 506420 -800 506532 480
rect 507602 -800 507714 480
rect 508784 -800 508896 480
rect 509966 -800 510078 480
rect 511148 -800 511260 480
rect 512330 -800 512442 480
rect 513512 -800 513624 480
rect 514694 -800 514806 480
rect 515876 -800 515988 480
rect 517058 -800 517170 480
rect 518240 -800 518352 480
rect 519422 -800 519534 480
rect 520604 -800 520716 480
rect 521786 -800 521898 480
rect 522968 -800 523080 480
rect 524150 -800 524262 480
rect 525332 -800 525444 480
rect 526514 -800 526626 480
rect 527696 -800 527808 480
rect 528878 -800 528990 480
rect 530060 -800 530172 480
rect 531242 -800 531354 480
rect 532424 -800 532536 480
rect 533606 -800 533718 480
rect 534788 -800 534900 480
rect 535970 -800 536082 480
rect 537152 -800 537264 480
rect 538334 -800 538446 480
rect 539516 -800 539628 480
rect 540698 -800 540810 480
rect 541880 -800 541992 480
rect 543062 -800 543174 480
rect 544244 -800 544356 480
rect 545426 -800 545538 480
rect 546608 -800 546720 480
rect 547790 -800 547902 480
rect 548972 -800 549084 480
rect 550154 -800 550266 480
rect 551336 -800 551448 480
rect 552518 -800 552630 480
rect 553700 -800 553812 480
rect 554882 -800 554994 480
rect 556064 -800 556176 480
rect 557246 -800 557358 480
rect 558428 -800 558540 480
rect 559610 -800 559722 480
rect 560792 -800 560904 480
rect 561974 -800 562086 480
rect 563156 -800 563268 480
rect 564338 -800 564450 480
rect 565520 -800 565632 480
rect 566702 -800 566814 480
rect 567884 -800 567996 480
rect 569066 -800 569178 480
rect 570248 -800 570360 480
rect 571430 -800 571542 480
rect 572612 -800 572724 480
rect 573794 -800 573906 480
rect 574976 -800 575088 480
rect 576158 -800 576270 480
rect 577340 -800 577452 480
rect 578522 -800 578634 480
rect 579704 -800 579816 480
rect 580886 -800 580998 480
rect 582068 -800 582180 480
rect 583250 -800 583362 480
<< via2 >>
rect 119008 695156 119292 695430
rect 120660 694918 121252 695446
rect 121760 694918 122352 695446
rect 122860 694918 123452 695446
rect 123960 694918 124552 695446
rect 126230 695110 126562 695464
rect 415392 691208 415494 691316
rect 415752 691208 415854 691316
rect 415392 690968 415494 691076
rect 415752 690968 415854 691076
rect 467296 691308 467398 691416
rect 467656 691308 467758 691416
rect 467296 691068 467398 691176
rect 467656 691068 467758 691176
rect 569260 691308 569362 691416
rect 569620 691308 569722 691416
rect 569260 691068 569362 691176
rect 569620 691068 569722 691176
rect 571002 689284 571242 689592
rect 571002 688684 571242 688992
rect 413812 688212 413996 688376
rect 414212 688212 414396 688376
rect 67008 687156 67292 687430
rect 413812 687812 413996 687976
rect 414212 687812 414396 687976
rect 68660 686918 69252 687446
rect 69760 686918 70352 687446
rect 70860 686918 71452 687446
rect 71960 686918 72552 687446
rect 74230 687110 74562 687464
rect 413812 687412 413996 687576
rect 414212 687412 414396 687576
rect 413812 687012 413996 687176
rect 414212 687012 414396 687176
rect 416212 688212 416278 688376
rect 416278 688212 416396 688376
rect 416612 688212 416796 688376
rect 416212 687812 416278 687976
rect 416278 687812 416396 687976
rect 416612 687812 416796 687976
rect 416212 687412 416278 687576
rect 416278 687412 416396 687576
rect 416612 687412 416796 687576
rect 416212 687012 416278 687176
rect 416278 687012 416396 687176
rect 416622 687012 416806 687176
rect 465812 688212 465996 688376
rect 466212 688212 466396 688376
rect 465812 687812 465996 687976
rect 466212 687812 466396 687976
rect 465812 687412 465996 687576
rect 466212 687412 466396 687576
rect 465812 687012 465996 687176
rect 466212 687012 466396 687176
rect 468212 688212 468396 688376
rect 468612 688212 468796 688376
rect 468212 687812 468396 687976
rect 468612 687812 468796 687976
rect 468212 687412 468396 687576
rect 468612 687412 468796 687576
rect 468212 687012 468396 687176
rect 468622 687012 468806 687176
rect 568212 688212 568396 688376
rect 568612 688212 568796 688376
rect 568212 687812 568396 687976
rect 568612 687812 568796 687976
rect 568212 687412 568396 687576
rect 568612 687412 568796 687576
rect 568212 687012 568396 687176
rect 568622 687012 568806 687176
rect 571002 688084 571242 688392
rect 571002 687484 571242 687792
rect 571002 686884 571242 687192
rect 571002 686284 571242 686592
rect 571002 685684 571242 685992
rect 415606 685408 415708 685516
rect 415966 685408 416068 685516
rect 415606 685168 415708 685276
rect 415966 685168 416068 685276
rect 467190 685404 467292 685512
rect 467550 685404 467652 685512
rect 467190 685164 467292 685272
rect 467550 685164 467652 685272
rect 569256 683708 569260 683814
rect 569260 683708 569362 683814
rect 569362 683708 569620 683814
rect 569620 683708 569722 683814
rect 569256 683576 569722 683708
rect 569256 683468 569260 683576
rect 569260 683468 569362 683576
rect 569362 683468 569620 683576
rect 569620 683468 569722 683576
rect 569256 683466 569722 683468
rect 70580 674824 70682 674932
rect 70940 674824 71042 674932
rect 70580 674584 70682 674692
rect 70940 674584 71042 674692
rect 122568 674866 122670 674974
rect 122928 674866 123030 674974
rect 122568 674626 122670 674734
rect 122928 674626 123030 674734
rect 70008 673458 70292 673732
rect 71368 673402 71700 673756
rect 121808 673220 122092 673494
rect 123302 673110 123634 673464
rect 70570 672224 70672 672332
rect 70930 672224 71032 672332
rect 70570 671984 70672 672092
rect 70930 671984 71032 672092
rect 122558 672266 122660 672374
rect 122918 672266 123020 672374
rect 122558 672026 122660 672134
rect 122918 672026 123020 672134
rect 440252 593576 440354 593684
rect 440612 593576 440714 593684
rect 440252 593336 440354 593444
rect 440612 593336 440714 593444
rect 448600 593608 448702 593716
rect 448960 593608 449062 593716
rect 448600 593368 448702 593476
rect 448960 593368 449062 593476
rect 437812 591984 437996 592148
rect 438212 591984 438396 592148
rect 437812 591584 437996 591748
rect 438212 591584 438396 591748
rect 437812 591184 437996 591348
rect 438212 591184 438396 591348
rect 437812 590784 437996 590948
rect 438212 590784 438396 590948
rect 442412 592080 442596 592244
rect 442812 592080 442996 592244
rect 442412 591680 442596 591844
rect 442812 591680 442996 591844
rect 442412 591280 442596 591444
rect 442812 591280 442996 591444
rect 442412 590880 442596 591044
rect 442822 590880 443006 591044
rect 446212 591984 446396 592148
rect 446612 591984 446796 592148
rect 446212 591584 446396 591748
rect 446612 591584 446796 591748
rect 446212 591184 446396 591348
rect 446612 591184 446796 591348
rect 446212 590784 446396 590948
rect 446612 590784 446796 590948
rect 450812 592080 450996 592244
rect 451212 592080 451396 592244
rect 450812 591680 450996 591844
rect 451212 591680 451396 591844
rect 450812 591280 450996 591444
rect 451212 591280 451396 591444
rect 450812 590880 450996 591044
rect 451222 590880 451406 591044
rect 440260 590104 440362 590212
rect 440620 590104 440722 590212
rect 440260 589864 440362 589972
rect 440620 589864 440722 589972
rect 448588 590104 448690 590212
rect 448948 590104 449050 590212
rect 448588 589864 448690 589972
rect 448948 589864 449050 589972
rect 405560 588304 405868 588544
rect 406160 588304 406468 588544
rect 406760 588304 407068 588544
rect 407360 588304 407668 588544
rect 407960 588304 408268 588544
rect 408560 588304 408868 588544
rect 409160 588304 409468 588544
rect 405006 587640 405086 587696
rect 405126 587640 405206 587696
rect 405006 587540 405086 587596
rect 405126 587540 405206 587596
rect 409990 587640 410070 587696
rect 410110 587640 410190 587696
rect 409990 587540 410070 587596
rect 410110 587540 410190 587596
rect 405560 586104 405868 586344
rect 406160 586104 406468 586344
rect 406760 586104 407068 586344
rect 407360 586104 407668 586344
rect 407960 586104 408268 586344
rect 408560 586104 408868 586344
rect 409160 586104 409468 586344
rect 416472 585948 417092 586336
rect 438974 586180 441846 586394
rect 405006 585540 405086 585596
rect 405126 585540 405206 585596
rect 405006 585440 405086 585496
rect 405126 585440 405206 585496
rect 409998 585540 410078 585596
rect 410118 585540 410198 585596
rect 409998 585440 410078 585496
rect 410118 585440 410198 585496
rect 416474 584828 417094 585216
rect 447368 584840 450242 585042
rect 405622 580628 406400 581174
rect 406822 580628 407600 581174
rect 408022 580628 408800 581174
rect 409222 580628 410000 581174
<< metal3 >>
rect 16194 702300 21194 704800
rect 68194 702928 73194 704800
rect 120194 703294 125194 704800
rect 68150 691494 73222 702928
rect 120124 695548 125196 703294
rect 165594 700170 170596 704800
rect 170894 702714 173094 704800
rect 165578 698240 170596 700170
rect 170854 702300 173094 702714
rect 173394 703810 175594 704800
rect 173394 702300 175744 703810
rect 175896 702300 180896 704800
rect 217294 702300 222294 704800
rect 222594 703328 224794 704800
rect 222500 702300 224794 703328
rect 225094 702300 227294 704800
rect 227594 702300 232594 704800
rect 318994 702300 323994 704800
rect 324294 702300 326494 704800
rect 326794 702300 328994 704800
rect 329294 702300 334294 704800
rect 413394 703906 418394 704800
rect 413390 702300 418394 703906
rect 465394 702880 470394 704800
rect 510594 702892 515394 704800
rect 118982 695430 119314 695454
rect 118982 695156 119008 695430
rect 119292 695156 119314 695430
rect 118982 695134 119314 695156
rect 120124 695446 125194 695548
rect 120124 694918 120660 695446
rect 121252 694918 121760 695446
rect 122352 694918 122860 695446
rect 123452 694918 123960 695446
rect 124552 695442 125194 695446
rect 126152 695464 126622 695524
rect 124552 694918 125196 695442
rect 126152 695110 126230 695464
rect 126562 695110 126622 695464
rect 126152 695052 126622 695110
rect 120124 693214 125196 694918
rect 119960 692034 125224 693214
rect 170854 692700 173082 702300
rect 170832 692140 173082 692700
rect 68096 691136 73222 691494
rect 68096 689728 73170 691136
rect 68096 687716 73196 689728
rect 68096 687454 73194 687716
rect 74152 687464 74622 687524
rect 66982 687430 67314 687454
rect 66982 687156 67008 687430
rect 67292 687156 67314 687430
rect 66982 687134 67314 687156
rect 68096 687446 73512 687454
rect 68096 686918 68660 687446
rect 69252 686918 69760 687446
rect 70352 686918 70860 687446
rect 71452 686918 71960 687446
rect 72552 687156 73512 687446
rect 72552 686919 73194 687156
rect 74152 687110 74230 687464
rect 74562 687110 74622 687464
rect 74152 687052 74622 687110
rect 72552 686918 73196 686919
rect 68096 685364 73196 686918
rect -800 680242 1700 685242
rect 68096 683432 73170 685364
rect 68096 683228 73222 683432
rect 68150 676930 73222 683228
rect 68130 674932 73246 676930
rect 68130 674824 70580 674932
rect 70682 674824 70940 674932
rect 71042 674824 73246 674932
rect 68130 674692 73246 674824
rect 68130 674584 70580 674692
rect 70682 674584 70940 674692
rect 71042 674584 73246 674692
rect 68130 674274 73246 674584
rect 120124 674974 125196 692034
rect 120124 674866 122568 674974
rect 122670 674866 122928 674974
rect 123030 674866 125196 674974
rect 120124 674734 125196 674866
rect 120124 674626 122568 674734
rect 122670 674626 122928 674734
rect 123030 674626 125196 674734
rect 120124 674080 125196 674626
rect 170832 674608 173060 692140
rect 71290 673756 71760 673816
rect 69982 673732 70314 673756
rect 69982 673458 70008 673732
rect 70292 673458 70314 673732
rect 69982 673436 70314 673458
rect 71290 673402 71368 673756
rect 71700 673402 71760 673756
rect 71290 673344 71760 673402
rect 121782 673494 122114 673518
rect 121782 673220 121808 673494
rect 122092 673220 122114 673494
rect 121782 673198 122114 673220
rect 123224 673464 123694 673524
rect 123224 673110 123302 673464
rect 123634 673110 123694 673464
rect 123224 673052 123694 673110
rect 68120 672332 73236 672874
rect 68120 672224 70570 672332
rect 70672 672224 70930 672332
rect 71032 672224 73236 672332
rect 68120 672092 73236 672224
rect 68120 671984 70570 672092
rect 70672 671984 70930 672092
rect 71032 671984 73236 672092
rect 68120 670218 73236 671984
rect 120124 672660 122044 672662
rect 123754 672660 125196 672662
rect 120124 672374 125196 672660
rect 170832 672644 173078 674608
rect 120124 672266 122558 672374
rect 122660 672266 122918 672374
rect 123020 672266 125196 672374
rect 120124 672134 125196 672266
rect 120124 672026 122558 672134
rect 122660 672026 122918 672134
rect 123020 672026 125196 672134
rect -800 643842 1660 648642
rect -800 633842 1660 638642
rect 68150 619820 73222 670218
rect 68150 618130 73250 619820
rect 120124 619052 125196 672026
rect 170720 664214 173078 672644
rect 170584 663610 173078 664214
rect 170584 656290 171186 663610
rect 172478 662146 173078 663610
rect 172478 656290 172824 662146
rect 170584 655688 172824 656290
rect 173464 644306 175744 702300
rect 222500 664812 224720 702300
rect 222260 664238 224752 664812
rect 222260 656624 222764 664238
rect 224356 656624 224752 664238
rect 222260 656278 224752 656624
rect 225202 657302 227234 702300
rect 413390 691862 418372 702300
rect 465390 697902 470394 702880
rect 465384 693606 470396 697902
rect 510580 696352 515412 702892
rect 520594 702688 525394 704800
rect 566594 702718 571594 704800
rect 520592 696352 525424 702688
rect 566588 700578 571618 702718
rect 529252 698920 531808 698936
rect 566584 698928 571618 700578
rect 534454 698920 562532 698928
rect 529252 698820 562532 698920
rect 529252 696842 564174 698820
rect 529252 696792 531808 696842
rect 534454 696828 564174 696842
rect 566536 696828 571618 698928
rect 510580 695166 525452 696352
rect 465384 693418 470416 693606
rect 465390 693184 470416 693418
rect 465392 692464 470416 693184
rect 465390 691986 470416 692464
rect 413348 691316 418396 691862
rect 413348 691208 415392 691316
rect 415494 691208 415752 691316
rect 415854 691208 418396 691316
rect 413348 691076 418396 691208
rect 413348 690968 415392 691076
rect 415494 690968 415752 691076
rect 415854 690968 418396 691076
rect 413348 689420 418396 690968
rect 465356 691562 470416 691986
rect 510494 691578 525452 695166
rect 465356 691416 470418 691562
rect 465356 691308 467296 691416
rect 467398 691308 467656 691416
rect 467758 691308 470418 691416
rect 465356 691176 470418 691308
rect 465356 691068 467296 691176
rect 467398 691068 467656 691176
rect 467758 691068 470418 691176
rect 465356 690870 470418 691068
rect 465356 689904 470396 690870
rect 413730 688376 414462 688608
rect 413730 688212 413812 688376
rect 413996 688212 414212 688376
rect 414396 688212 414462 688376
rect 413730 687976 414462 688212
rect 413730 687812 413812 687976
rect 413996 687812 414212 687976
rect 414396 687812 414462 687976
rect 413730 687576 414462 687812
rect 413730 687412 413812 687576
rect 413996 687412 414212 687576
rect 414396 687412 414462 687576
rect 413730 687176 414462 687412
rect 413730 687012 413812 687176
rect 413996 687012 414212 687176
rect 414396 687012 414462 687176
rect 413730 686944 414462 687012
rect 416130 688376 416866 688598
rect 416130 688212 416212 688376
rect 416396 688212 416612 688376
rect 416796 688212 416866 688376
rect 416130 687976 416866 688212
rect 416130 687812 416212 687976
rect 416396 687812 416612 687976
rect 416796 687812 416866 687976
rect 416130 687576 416866 687812
rect 416130 687412 416212 687576
rect 416396 687412 416612 687576
rect 416796 687412 416866 687576
rect 416130 687176 416866 687412
rect 416130 687012 416212 687176
rect 416396 687012 416622 687176
rect 416806 687012 416866 687176
rect 416130 686944 416866 687012
rect 465730 688376 466466 688608
rect 465730 688212 465812 688376
rect 465996 688212 466212 688376
rect 466396 688212 466466 688376
rect 465730 687976 466466 688212
rect 465730 687812 465812 687976
rect 465996 687812 466212 687976
rect 466396 687812 466466 687976
rect 465730 687576 466466 687812
rect 465730 687412 465812 687576
rect 465996 687412 466212 687576
rect 466396 687412 466466 687576
rect 465730 687176 466466 687412
rect 465730 687012 465812 687176
rect 465996 687012 466212 687176
rect 466396 687012 466466 687176
rect 465730 686944 466466 687012
rect 468130 688376 468866 688598
rect 468130 688212 468212 688376
rect 468396 688212 468612 688376
rect 468796 688212 468866 688376
rect 468130 687976 468866 688212
rect 468130 687812 468212 687976
rect 468396 687812 468612 687976
rect 468796 687812 468866 687976
rect 468130 687576 468866 687812
rect 468130 687412 468212 687576
rect 468396 687412 468612 687576
rect 468796 687412 468866 687576
rect 468130 687176 468866 687412
rect 468130 687012 468212 687176
rect 468396 687012 468622 687176
rect 468806 687012 468866 687176
rect 468130 686944 468866 687012
rect 510494 686746 512924 691578
rect 517294 686746 519782 691578
rect 524152 687904 525452 691578
rect 524152 686746 525424 687904
rect 413382 685516 418382 685878
rect 466946 685578 467272 685580
rect 466650 685576 468836 685578
rect 465390 685546 470376 685576
rect 413382 685408 415606 685516
rect 415708 685408 415966 685516
rect 416068 685408 418382 685516
rect 413382 685276 418382 685408
rect 413382 685168 415606 685276
rect 415708 685168 415966 685276
rect 416068 685168 418382 685276
rect 413382 685074 418382 685168
rect 465318 685512 470376 685546
rect 465318 685404 467190 685512
rect 467292 685404 467550 685512
rect 467652 685404 470376 685512
rect 465318 685272 470376 685404
rect 465318 685164 467190 685272
rect 467292 685164 467550 685272
rect 467652 685164 470376 685272
rect 413388 684800 418376 685074
rect 465318 684800 470376 685164
rect 413390 672446 418372 684800
rect 465318 684084 470372 684800
rect 510494 684518 525424 686746
rect 465318 683036 470370 684084
rect 465318 682080 470394 683036
rect 465390 672488 470394 682080
rect 426718 672486 433774 672488
rect 426718 672446 441922 672486
rect 413390 667906 441922 672446
rect 438918 659596 441922 667906
rect 447300 667914 470394 672488
rect 447300 667900 451926 667914
rect 447318 661028 450322 667900
rect 465390 667864 470394 667914
rect 529252 669536 531138 696792
rect 534982 691808 543812 693940
rect 529252 667346 531270 669536
rect 438868 658800 441950 659596
rect 447318 659006 450330 661028
rect 438868 658322 441984 658800
rect 225202 656220 227256 657302
rect 173466 641340 175738 644306
rect 216098 641350 221908 641414
rect 225206 641350 227256 656220
rect 438908 652464 441984 658322
rect 447312 652670 450388 659006
rect 438924 651142 441968 652464
rect 438918 650114 441968 651142
rect 447316 651142 450320 652670
rect 227664 641350 238982 641414
rect 163350 641316 170068 641340
rect 160032 641306 170068 641316
rect 173362 641316 179734 641340
rect 216098 641316 238982 641350
rect 351700 641316 362636 641330
rect 160032 641300 172954 641306
rect 173362 641300 362636 641316
rect 160032 639526 362636 641300
rect 160032 633438 354208 639526
rect 360382 633438 362636 639526
rect 160032 631774 362636 633438
rect 160032 631742 167582 631774
rect 177012 631742 362636 631774
rect 216098 631660 238982 631742
rect 351700 631718 362636 631742
rect 68154 613838 73250 618130
rect 68150 612936 73250 613838
rect 68150 593482 73222 612936
rect 119910 611580 125354 619052
rect 67942 585606 73258 593482
rect 119960 587712 125224 611580
rect 438918 593684 441922 650114
rect 447316 649884 450322 651142
rect 438918 593576 440252 593684
rect 440354 593576 440612 593684
rect 440714 593576 441922 593684
rect 438918 593444 441922 593576
rect 438918 593336 440252 593444
rect 440354 593336 440612 593444
rect 440714 593336 441922 593444
rect 438918 592640 441922 593336
rect 447318 593716 450322 649884
rect 529258 646566 531270 667346
rect 535058 646566 536962 691808
rect 542138 667672 543812 691808
rect 548912 691712 557742 693844
rect 529258 645074 536962 646566
rect 542034 646524 543894 667672
rect 548972 646524 550582 691712
rect 556032 647396 557702 691712
rect 562262 684168 564174 696828
rect 566584 696820 571618 696828
rect 566584 693830 571614 696820
rect 566562 691712 571632 693830
rect 566562 691416 571616 691712
rect 566562 691308 569260 691416
rect 569362 691308 569620 691416
rect 569722 691308 571616 691416
rect 566562 691176 571616 691308
rect 566562 691068 569260 691176
rect 569362 691068 569620 691176
rect 569722 691068 571616 691176
rect 566562 690650 571616 691068
rect 570922 689592 571352 689764
rect 570922 689284 571002 689592
rect 571242 689284 571352 689592
rect 570922 688992 571352 689284
rect 570922 688684 571002 688992
rect 571242 688684 571352 688992
rect 568130 688376 568866 688598
rect 568130 688212 568212 688376
rect 568396 688212 568612 688376
rect 568796 688212 568866 688376
rect 568130 687976 568866 688212
rect 568130 687812 568212 687976
rect 568396 687812 568612 687976
rect 568796 687812 568866 687976
rect 568130 687576 568866 687812
rect 568130 687412 568212 687576
rect 568396 687412 568612 687576
rect 568796 687412 568866 687576
rect 568130 687176 568866 687412
rect 568130 687012 568212 687176
rect 568396 687012 568622 687176
rect 568806 687012 568866 687176
rect 568130 686944 568866 687012
rect 570922 688392 571352 688684
rect 570922 688084 571002 688392
rect 571242 688084 571352 688392
rect 570922 687792 571352 688084
rect 570922 687484 571002 687792
rect 571242 687484 571352 687792
rect 570922 687192 571352 687484
rect 570922 686884 571002 687192
rect 571242 686884 571352 687192
rect 570922 686592 571352 686884
rect 570922 686284 571002 686592
rect 571242 686284 571352 686592
rect 570922 685992 571352 686284
rect 570922 685684 571002 685992
rect 571242 685684 571352 685992
rect 570922 685072 571352 685684
rect 562262 683814 570108 684168
rect 562262 683466 569256 683814
rect 569722 683466 570108 683814
rect 562262 683252 570108 683466
rect 562296 681638 570108 683252
rect 572674 683000 577382 683012
rect 572674 682984 583000 683000
rect 572674 677996 584800 682984
rect 572674 676228 577382 677996
rect 582300 677984 584800 677996
rect 562824 675840 577382 676228
rect 562780 671002 577382 675840
rect 562780 670958 576172 671002
rect 562780 668898 564676 670958
rect 562780 660762 564594 668898
rect 562862 647396 564532 660762
rect 556032 647266 564600 647396
rect 542034 645242 550582 646524
rect 556056 645904 564600 647266
rect 529258 645056 531270 645074
rect 535058 644996 536962 645074
rect 542038 645032 550582 645242
rect 548972 644982 550582 645032
rect 565206 644596 576142 646006
rect 565206 644584 583128 644596
rect 565206 644560 584800 644584
rect 565206 641590 567706 644560
rect 564368 639756 567706 641590
rect 573760 639812 584800 644560
rect 573760 639756 576142 639812
rect 582340 639784 584800 639812
rect 564368 634590 576142 639756
rect 564368 634584 583082 634590
rect 564368 634562 584800 634584
rect 564368 632060 567668 634562
rect 565206 629758 567668 632060
rect 573722 629784 584800 634562
rect 573722 629758 576142 629784
rect 565206 627532 576142 629758
rect 447318 593608 448600 593716
rect 448702 593608 448960 593716
rect 449062 593608 450322 593716
rect 447318 593476 450322 593608
rect 447318 593368 448600 593476
rect 448702 593368 448960 593476
rect 449062 593368 450322 593476
rect 438920 592518 441916 592640
rect 447318 592624 450322 593368
rect 437730 592148 438466 592380
rect 437730 591984 437812 592148
rect 437996 591984 438212 592148
rect 438396 591984 438466 592148
rect 437730 591748 438466 591984
rect 437730 591584 437812 591748
rect 437996 591584 438212 591748
rect 438396 591584 438466 591748
rect 437730 591348 438466 591584
rect 437730 591184 437812 591348
rect 437996 591184 438212 591348
rect 438396 591184 438466 591348
rect 437730 590948 438466 591184
rect 437730 590784 437812 590948
rect 437996 590784 438212 590948
rect 438396 590784 438466 590948
rect 442330 592244 443066 592420
rect 442330 592080 442412 592244
rect 442596 592080 442812 592244
rect 442996 592080 443066 592244
rect 442330 591844 443066 592080
rect 442330 591680 442412 591844
rect 442596 591680 442812 591844
rect 442996 591680 443066 591844
rect 442330 591444 443066 591680
rect 442330 591280 442412 591444
rect 442596 591280 442812 591444
rect 442996 591280 443066 591444
rect 442330 591044 443066 591280
rect 442330 590880 442412 591044
rect 442596 590880 442822 591044
rect 443006 590880 443066 591044
rect 442330 590812 443066 590880
rect 446130 592148 446866 592380
rect 446130 591984 446212 592148
rect 446396 591984 446612 592148
rect 446796 591984 446866 592148
rect 446130 591748 446866 591984
rect 446130 591584 446212 591748
rect 446396 591584 446612 591748
rect 446796 591584 446866 591748
rect 446130 591348 446866 591584
rect 446130 591184 446212 591348
rect 446396 591184 446612 591348
rect 446796 591184 446866 591348
rect 446130 590948 446866 591184
rect 437730 590716 438466 590784
rect 446130 590784 446212 590948
rect 446396 590784 446612 590948
rect 446796 590784 446866 590948
rect 450730 592244 451466 592420
rect 450730 592080 450812 592244
rect 450996 592080 451212 592244
rect 451396 592080 451466 592244
rect 450730 591844 451466 592080
rect 450730 591680 450812 591844
rect 450996 591680 451212 591844
rect 451396 591680 451466 591844
rect 450730 591444 451466 591680
rect 450730 591280 450812 591444
rect 450996 591280 451212 591444
rect 451396 591280 451466 591444
rect 450730 591044 451466 591280
rect 450730 590880 450812 591044
rect 450996 590880 451222 591044
rect 451406 590880 451466 591044
rect 450730 590812 451466 590880
rect 446130 590716 446866 590784
rect 439822 590556 441246 590562
rect 448222 590556 449646 590562
rect 438918 590212 441922 590556
rect 438918 590104 440260 590212
rect 440362 590104 440620 590212
rect 440722 590104 441922 590212
rect 438918 589972 441922 590104
rect 438918 589864 440260 589972
rect 440362 589864 440620 589972
rect 440722 589864 441922 589972
rect 405388 588544 410080 588654
rect 405388 588304 405560 588544
rect 405868 588304 406160 588544
rect 406468 588304 406760 588544
rect 407068 588304 407360 588544
rect 407668 588304 407960 588544
rect 408268 588304 408560 588544
rect 408868 588304 409160 588544
rect 409468 588304 410080 588544
rect 405388 588224 410080 588304
rect 415556 587732 415682 587738
rect 225668 587714 233592 587722
rect 218102 587712 233592 587714
rect 404834 587712 405254 587728
rect 119960 587696 405254 587712
rect 409972 587710 411912 587714
rect 415556 587712 417000 587732
rect 412282 587710 417000 587712
rect 409972 587706 421224 587710
rect 119960 587640 405006 587696
rect 405086 587640 405126 587696
rect 405206 587640 405254 587696
rect 119960 587596 405254 587640
rect 119960 587540 405006 587596
rect 405086 587540 405126 587596
rect 405206 587540 405254 587596
rect 119960 587528 405254 587540
rect 119960 587522 226026 587528
rect 119960 587518 203610 587522
rect 210580 587520 226026 587522
rect 210580 587518 218504 587520
rect 230148 587518 405254 587528
rect 119960 587514 129408 587518
rect 404286 587516 405254 587518
rect 119960 587492 125224 587514
rect 404834 587472 405254 587516
rect 409966 587700 421224 587706
rect 409966 587696 421478 587700
rect 409966 587640 409990 587696
rect 410070 587640 410110 587696
rect 410190 587640 421478 587696
rect 409966 587596 421478 587640
rect 409966 587540 409990 587596
rect 410070 587540 410110 587596
rect 410190 587540 421478 587596
rect 409966 587518 421478 587540
rect 409966 587512 412420 587518
rect 415568 587516 421478 587518
rect 415568 587512 417000 587516
rect 409968 587510 410212 587512
rect 411726 587510 412420 587512
rect 421078 586934 421478 587516
rect 405388 586344 410080 586454
rect 405388 586104 405560 586344
rect 405868 586104 406160 586344
rect 406468 586104 406760 586344
rect 407068 586104 407360 586344
rect 407668 586104 407960 586344
rect 408268 586104 408560 586344
rect 408868 586104 409160 586344
rect 409468 586104 410080 586344
rect 405388 586024 410080 586104
rect 416354 586336 417192 586444
rect 438918 586394 441922 589864
rect 447318 590212 450322 590556
rect 447318 590104 448588 590212
rect 448690 590104 448948 590212
rect 449050 590104 450322 590212
rect 447318 589972 450322 590104
rect 447318 589864 448588 589972
rect 448690 589864 448948 589972
rect 449050 589864 450322 589972
rect 447318 586662 450322 589864
rect 583520 589472 584800 589584
rect 583520 588290 584800 588402
rect 583520 587108 584800 587220
rect 447316 586398 450322 586662
rect 438918 586356 438974 586394
rect 416354 585948 416472 586336
rect 417092 585948 417192 586336
rect 438908 586180 438974 586356
rect 441846 586356 441922 586394
rect 441846 586180 441924 586356
rect 438908 586102 441924 586180
rect 447312 586048 450322 586398
rect 416354 585850 417192 585948
rect 416094 585606 417324 585612
rect 67942 585604 218504 585606
rect 230148 585604 405258 585606
rect 67942 585596 405258 585604
rect 67942 585540 405006 585596
rect 405086 585540 405126 585596
rect 405206 585540 405258 585596
rect 67942 585496 405258 585540
rect 67942 585440 405006 585496
rect 405086 585440 405126 585496
rect 405206 585440 405258 585496
rect 67942 585412 405258 585440
rect 409974 585596 417324 585606
rect 409974 585540 409998 585596
rect 410078 585540 410118 585596
rect 410198 585540 417324 585596
rect 409974 585496 417324 585540
rect 409974 585440 409998 585496
rect 410078 585440 410118 585496
rect 410198 585440 417324 585496
rect 409974 585416 417324 585440
rect 409974 585412 416016 585416
rect 416354 585414 417186 585416
rect 447316 585414 450318 586048
rect 583520 585926 584800 586038
rect 67942 585282 73258 585412
rect 218288 585410 230804 585412
rect 404984 585410 405258 585412
rect 409976 585410 410220 585412
rect 415798 585408 416016 585412
rect 416356 585216 417188 585316
rect 416356 584828 416474 585216
rect 417094 584828 417188 585216
rect 416356 584730 417188 584828
rect 447312 585258 450318 585414
rect 447312 585042 450316 585258
rect 447312 584840 447368 585042
rect 450242 584840 450316 585042
rect 447312 584780 450316 584840
rect 583520 584744 584800 584856
rect 583520 583562 584800 583674
rect 405234 581174 410146 581588
rect 405234 580628 405622 581174
rect 406400 580628 406822 581174
rect 407600 580628 408022 581174
rect 408800 580628 409222 581174
rect 410000 580628 410146 581174
rect 405234 580232 410146 580628
rect -800 559442 1660 564242
rect -800 549442 1660 554242
rect 582340 550562 584800 555362
rect 582340 540562 584800 545362
rect -800 511530 480 511642
rect -800 510348 480 510460
rect -800 509166 480 509278
rect -800 507984 480 508096
rect -800 506802 480 506914
rect -800 505620 480 505732
rect 583520 500050 584800 500162
rect 583520 498868 584800 498980
rect 583520 497686 584800 497798
rect 583520 496504 584800 496616
rect 583520 495322 584800 495434
rect 583520 494140 584800 494252
rect -800 468308 480 468420
rect -800 467126 480 467238
rect -800 465944 480 466056
rect -800 464762 480 464874
rect -800 463580 480 463692
rect -800 462398 480 462510
rect 583520 455628 584800 455740
rect 583520 454446 584800 454558
rect 583520 453264 584800 453376
rect 583520 452082 584800 452194
rect 583520 450900 584800 451012
rect 583520 449718 584800 449830
rect -800 425086 480 425198
rect -800 423904 480 424016
rect -800 422722 480 422834
rect -800 421540 480 421652
rect -800 420358 480 420470
rect -800 419176 480 419288
rect 583520 411206 584800 411318
rect 583520 410024 584800 410136
rect 583520 408842 584800 408954
rect 583520 407660 584800 407772
rect 583520 406478 584800 406590
rect 583520 405296 584800 405408
rect -800 381864 480 381976
rect -800 380682 480 380794
rect -800 379500 480 379612
rect -800 378318 480 378430
rect -800 377136 480 377248
rect -800 375954 480 376066
rect 583520 364784 584800 364896
rect 583520 363602 584800 363714
rect 583520 362420 584800 362532
rect 583520 361238 584800 361350
rect 583520 360056 584800 360168
rect 583520 358874 584800 358986
rect -800 338642 480 338754
rect -800 337460 480 337572
rect -800 336278 480 336390
rect -800 335096 480 335208
rect -800 333914 480 334026
rect -800 332732 480 332844
rect 583520 319562 584800 319674
rect 583520 318380 584800 318492
rect 583520 317198 584800 317310
rect 583520 316016 584800 316128
rect 583520 314834 584800 314946
rect 583520 313652 584800 313764
rect -800 295420 480 295532
rect -800 294238 480 294350
rect -800 293056 480 293168
rect -800 291874 480 291986
rect -800 290692 480 290804
rect -800 289510 480 289622
rect 583520 275140 584800 275252
rect 583520 273958 584800 274070
rect 583520 272776 584800 272888
rect 583520 271594 584800 271706
rect 583520 270412 584800 270524
rect 583520 269230 584800 269342
rect -800 252398 480 252510
rect -800 251216 480 251328
rect -800 250034 480 250146
rect -800 248852 480 248964
rect -800 247670 480 247782
rect -800 246488 480 246600
rect 582340 235230 584800 240030
rect 582340 225230 584800 230030
rect -800 214888 1660 219688
rect -800 204888 1660 209688
rect 582188 196230 582876 196238
rect 582188 191430 584800 196230
rect 582188 191424 582876 191430
rect 582340 186224 584800 186230
rect 582188 181430 584800 186224
rect 582188 181410 582678 181430
rect -800 172888 1660 177688
rect -800 162888 1660 167688
rect 582340 151538 584800 151630
rect 581994 146830 584800 151538
rect 581994 146778 583364 146830
rect 581994 141630 583088 141672
rect 581994 136912 584800 141630
rect 582340 136830 584800 136912
rect -800 124776 480 124888
rect -800 123594 480 123706
rect -800 122412 480 122524
rect -800 121230 480 121342
rect -800 120048 480 120160
rect -800 118866 480 118978
rect 583520 95118 584800 95230
rect 583520 93936 584800 94048
rect 583520 92754 584800 92866
rect 583520 91572 584800 91684
rect -800 81554 480 81666
rect -800 80372 480 80484
rect -800 79190 480 79302
rect -800 78008 480 78120
rect -800 76826 480 76938
rect -800 75644 480 75756
rect 583520 50460 584800 50572
rect 583520 49278 584800 49390
rect 583520 48096 584800 48208
rect 583520 46914 584800 47026
rect -800 38332 480 38444
rect -800 37150 480 37262
rect -800 35968 480 36080
rect -800 34786 480 34898
rect -800 33604 480 33716
rect -800 32422 480 32534
rect 583520 24002 584800 24114
rect 583520 22820 584800 22932
rect 583520 21638 584800 21750
rect 583520 20456 584800 20568
rect 583520 19274 584800 19386
rect 583520 18092 584800 18204
rect -800 16910 480 17022
rect 583520 16910 584800 17022
rect -800 15728 480 15840
rect 583520 15728 584800 15840
rect -800 14546 480 14658
rect 583520 14546 584800 14658
rect -800 13364 480 13476
rect 583520 13364 584800 13476
rect -800 12182 480 12294
rect 583520 12182 584800 12294
rect -800 11000 480 11112
rect 583520 11000 584800 11112
rect -800 9818 480 9930
rect 583520 9818 584800 9930
rect -800 8636 480 8748
rect 583520 8636 584800 8748
rect -800 7454 480 7566
rect 583520 7454 584800 7566
rect -800 6272 480 6384
rect 583520 6272 584800 6384
rect -800 5090 480 5202
rect 583520 5090 584800 5202
rect -800 3908 480 4020
rect 583520 3908 584800 4020
rect -800 2726 480 2838
rect 583520 2726 584800 2838
rect -800 1544 480 1656
rect 583520 1544 584800 1656
<< via3 >>
rect 119008 695156 119292 695430
rect 126230 695110 126562 695464
rect 67008 687156 67292 687430
rect 74230 687110 74562 687464
rect 70008 673458 70292 673732
rect 71368 673402 71700 673756
rect 121808 673220 122092 673494
rect 123302 673110 123634 673464
rect 171186 656290 172478 663610
rect 222764 656624 224356 664238
rect 413812 688212 413996 688376
rect 414212 688212 414396 688376
rect 413812 687812 413996 687976
rect 414212 687812 414396 687976
rect 413812 687412 413996 687576
rect 414212 687412 414396 687576
rect 413812 687012 413996 687176
rect 414212 687012 414396 687176
rect 416212 688212 416396 688376
rect 416612 688212 416796 688376
rect 416212 687812 416396 687976
rect 416612 687812 416796 687976
rect 416212 687412 416396 687576
rect 416612 687412 416796 687576
rect 416212 687012 416396 687176
rect 416622 687012 416806 687176
rect 465812 688212 465996 688376
rect 466212 688212 466396 688376
rect 465812 687812 465996 687976
rect 466212 687812 466396 687976
rect 465812 687412 465996 687576
rect 466212 687412 466396 687576
rect 465812 687012 465996 687176
rect 466212 687012 466396 687176
rect 468212 688212 468396 688376
rect 468612 688212 468796 688376
rect 468212 687812 468396 687976
rect 468612 687812 468796 687976
rect 468212 687412 468396 687576
rect 468612 687412 468796 687576
rect 468212 687012 468396 687176
rect 468622 687012 468806 687176
rect 512924 686746 517294 691578
rect 519782 686746 524152 691578
rect 354208 633438 360382 639526
rect 571002 689284 571242 689592
rect 571002 688684 571242 688992
rect 568212 688212 568396 688376
rect 568612 688212 568796 688376
rect 568212 687812 568396 687976
rect 568612 687812 568796 687976
rect 568212 687412 568396 687576
rect 568612 687412 568796 687576
rect 568212 687012 568396 687176
rect 568622 687012 568806 687176
rect 571002 688084 571242 688392
rect 571002 687484 571242 687792
rect 571002 686884 571242 687192
rect 571002 686284 571242 686592
rect 571002 685684 571242 685992
rect 567706 639756 573760 644560
rect 567668 629758 573722 634562
rect 437812 591984 437996 592148
rect 438212 591984 438396 592148
rect 437812 591584 437996 591748
rect 438212 591584 438396 591748
rect 437812 591184 437996 591348
rect 438212 591184 438396 591348
rect 437812 590784 437996 590948
rect 438212 590784 438396 590948
rect 442412 592080 442596 592244
rect 442812 592080 442996 592244
rect 442412 591680 442596 591844
rect 442812 591680 442996 591844
rect 442412 591280 442596 591444
rect 442812 591280 442996 591444
rect 442412 590880 442596 591044
rect 442822 590880 443006 591044
rect 446212 591984 446396 592148
rect 446612 591984 446796 592148
rect 446212 591584 446396 591748
rect 446612 591584 446796 591748
rect 446212 591184 446396 591348
rect 446612 591184 446796 591348
rect 446212 590784 446396 590948
rect 446612 590784 446796 590948
rect 450812 592080 450996 592244
rect 451212 592080 451396 592244
rect 450812 591680 450996 591844
rect 451212 591680 451396 591844
rect 450812 591280 450996 591444
rect 451212 591280 451396 591444
rect 450812 590880 450996 591044
rect 451222 590880 451406 591044
rect 405560 588304 405868 588544
rect 406160 588304 406468 588544
rect 406760 588304 407068 588544
rect 407360 588304 407668 588544
rect 407960 588304 408268 588544
rect 408560 588304 408868 588544
rect 409160 588304 409468 588544
rect 405560 586104 405868 586344
rect 406160 586104 406468 586344
rect 406760 586104 407068 586344
rect 407360 586104 407668 586344
rect 407960 586104 408268 586344
rect 408560 586104 408868 586344
rect 409160 586104 409468 586344
rect 416472 585948 417092 586336
rect 416474 584828 417094 585216
rect 405622 580628 406400 581174
rect 406822 580628 407600 581174
rect 408022 580628 408800 581174
rect 409222 580628 410000 581174
<< metal4 >>
rect 165594 700170 170596 704800
rect 175896 704714 180896 704800
rect 175894 702434 180896 704714
rect 217294 702970 222294 704800
rect 217294 702300 222298 702970
rect 227594 702926 232594 704800
rect 74154 687464 74702 687572
rect 86764 687466 98118 697602
rect 126154 695464 126702 695572
rect 118982 695430 119314 695454
rect 118982 695156 119008 695430
rect 119292 695156 119314 695430
rect 118982 695134 119314 695156
rect 126154 695110 126230 695464
rect 126562 695454 126702 695464
rect 136728 695456 148082 698648
rect 165578 698240 170596 700170
rect 217306 700998 222298 702300
rect 128578 695454 148082 695456
rect 126562 695134 148082 695454
rect 126562 695110 126698 695134
rect 128578 695132 148082 695134
rect 126154 694992 126698 695110
rect 66982 687430 67314 687454
rect 66982 687156 67008 687430
rect 67292 687156 67314 687430
rect 66982 687134 67314 687156
rect 74154 687110 74230 687464
rect 74562 687454 74702 687464
rect 75168 687454 98118 687466
rect 74562 687134 98118 687454
rect 74562 687110 74698 687134
rect 74154 686992 74698 687110
rect 86764 676416 98118 687134
rect 86766 674816 98118 676416
rect 136728 676412 148082 695132
rect 217306 684124 222336 700998
rect 170578 677212 175880 682686
rect 175818 677200 175880 677212
rect 180902 682660 187876 682686
rect 217280 682660 222336 684124
rect 227582 694624 232594 702926
rect 318994 702300 323994 704800
rect 329294 702300 334294 704800
rect 227582 682660 232548 694624
rect 402706 694056 464752 696958
rect 402738 688608 404890 694056
rect 463316 693774 464752 694056
rect 412670 688608 414760 688612
rect 463316 688610 464766 693774
rect 511622 691578 524816 694356
rect 402692 688376 414760 688608
rect 463308 688608 465444 688610
rect 416124 688598 416882 688604
rect 402692 688212 413812 688376
rect 413996 688212 414212 688376
rect 414396 688212 414760 688376
rect 402692 687976 414760 688212
rect 402692 687812 413812 687976
rect 413996 687812 414212 687976
rect 414396 687812 414760 687976
rect 402692 687576 414760 687812
rect 402692 687412 413812 687576
rect 413996 687412 414212 687576
rect 414396 687412 414760 687576
rect 402692 687176 414760 687412
rect 402692 687012 413812 687176
rect 413996 687012 414212 687176
rect 414396 687012 414760 687176
rect 402692 686948 414760 687012
rect 416120 688376 416882 688598
rect 416120 688212 416212 688376
rect 416396 688212 416612 688376
rect 416796 688212 416882 688376
rect 416120 688050 416882 688212
rect 416120 688042 416560 688050
rect 416120 687738 416166 688042
rect 416450 687746 416560 688042
rect 416844 687746 416882 688050
rect 416450 687738 416882 687746
rect 416120 687576 416882 687738
rect 416120 687412 416212 687576
rect 416396 687412 416612 687576
rect 416796 687412 416882 687576
rect 416120 687258 416882 687412
rect 416120 686962 416156 687258
rect 416484 687254 416882 687258
rect 416484 686962 416568 687254
rect 416120 686950 416568 686962
rect 416852 686950 416882 687254
rect 416120 686948 416882 686950
rect 180902 682658 191412 682660
rect 208250 682658 232548 682660
rect 180902 677212 191572 682658
rect 180902 677200 181542 677212
rect 185920 677168 191572 677212
rect 186724 676918 191572 677168
rect 204138 677168 232548 682658
rect 402730 681322 404890 686948
rect 412670 686942 414760 686948
rect 416124 686946 416882 686948
rect 463308 688376 466460 688608
rect 468124 688598 468882 688604
rect 463308 688212 465812 688376
rect 465996 688212 466212 688376
rect 466396 688212 466460 688376
rect 463308 687976 466460 688212
rect 463308 687812 465812 687976
rect 465996 687812 466212 687976
rect 466396 687812 466460 687976
rect 463308 687576 466460 687812
rect 463308 687412 465812 687576
rect 465996 687412 466212 687576
rect 466396 687412 466460 687576
rect 463308 687176 466460 687412
rect 463308 687012 465812 687176
rect 465996 687012 466212 687176
rect 466396 687012 466460 687176
rect 463308 686948 466460 687012
rect 468120 688376 468882 688598
rect 468120 688212 468212 688376
rect 468396 688212 468612 688376
rect 468796 688212 468882 688376
rect 468120 688050 468882 688212
rect 468120 688042 468560 688050
rect 468120 687738 468166 688042
rect 468450 687746 468560 688042
rect 468844 687746 468882 688050
rect 468450 687738 468882 687746
rect 468120 687576 468882 687738
rect 468120 687412 468212 687576
rect 468396 687412 468612 687576
rect 468796 687412 468882 687576
rect 468120 687258 468882 687412
rect 468120 686962 468156 687258
rect 468484 687254 468882 687258
rect 468484 686962 468568 687254
rect 468120 686950 468568 686962
rect 468852 686950 468882 687254
rect 468120 686948 468882 686950
rect 463308 686946 465444 686948
rect 468124 686946 468882 686948
rect 511622 686746 512924 691578
rect 517294 686746 519782 691578
rect 524152 686746 524816 691578
rect 571158 690202 575926 690212
rect 570574 689592 575926 690202
rect 570574 689284 571002 689592
rect 571242 689284 575926 689592
rect 570574 688992 575926 689284
rect 570574 688684 571002 688992
rect 571242 688684 575926 688992
rect 568124 688598 568882 688604
rect 568120 688376 568882 688598
rect 568120 688212 568212 688376
rect 568396 688212 568612 688376
rect 568796 688212 568882 688376
rect 568120 688050 568882 688212
rect 568120 688042 568560 688050
rect 568120 687738 568166 688042
rect 568450 687746 568560 688042
rect 568844 687746 568882 688050
rect 568450 687738 568882 687746
rect 568120 687576 568882 687738
rect 568120 687412 568212 687576
rect 568396 687412 568612 687576
rect 568796 687412 568882 687576
rect 568120 687258 568882 687412
rect 568120 686962 568156 687258
rect 568484 687254 568882 687258
rect 568484 686962 568568 687254
rect 568120 686950 568568 686962
rect 568852 686950 568882 687254
rect 568120 686948 568882 686950
rect 568124 686946 568882 686948
rect 570574 688392 575926 688684
rect 570574 688084 571002 688392
rect 571242 688084 575926 688392
rect 570574 687792 575926 688084
rect 570574 687484 571002 687792
rect 571242 687484 575926 687792
rect 570574 687192 575926 687484
rect 511622 684546 524816 686746
rect 570574 686884 571002 687192
rect 571242 686884 575926 687192
rect 570574 686592 575926 686884
rect 570574 686284 571002 686592
rect 571242 686284 575926 686592
rect 570574 685992 575926 686284
rect 570574 685684 571002 685992
rect 571242 685684 575926 685992
rect 570574 685480 575926 685684
rect 570574 683716 575942 685480
rect 204138 676918 209704 677168
rect 71292 673756 71840 673864
rect 78430 673758 81324 673770
rect 86764 673758 98118 674816
rect 69982 673732 70314 673756
rect 69982 673458 70008 673732
rect 70292 673458 70314 673732
rect 69982 673436 70314 673458
rect 71292 673402 71368 673756
rect 71700 673746 71840 673756
rect 75168 673746 98118 673758
rect 71700 673426 98118 673746
rect 71700 673402 71836 673426
rect 71292 673284 71836 673402
rect 86764 648996 98118 673426
rect 103262 673632 111234 675078
rect 136838 674412 148082 676412
rect 119710 673632 121470 673634
rect 103262 673494 122298 673632
rect 103262 673220 121808 673494
rect 122092 673220 122298 673494
rect 103262 673068 122298 673220
rect 123226 673464 123774 673572
rect 123226 673110 123302 673464
rect 123634 673454 123774 673464
rect 136728 673456 148082 674412
rect 128578 673454 148082 673456
rect 123634 673134 148082 673454
rect 123634 673110 123770 673134
rect 128578 673132 148082 673134
rect 103262 661186 111234 673068
rect 123226 672992 123770 673110
rect 99488 655198 111234 661186
rect 99464 654946 111234 655198
rect 99464 653892 111288 654946
rect 136728 650176 148082 673132
rect 222268 664238 224752 664696
rect 170584 663610 172824 664214
rect 170584 656290 171186 663610
rect 172478 661626 172824 663610
rect 222268 661626 222764 664238
rect 172478 661560 185306 661626
rect 213460 661560 222764 661626
rect 172478 658966 222764 661560
rect 172478 656290 172824 658966
rect 181400 658866 215482 658966
rect 170584 655688 172824 656290
rect 222268 656624 222764 658966
rect 224356 656624 224752 664238
rect 222268 656278 224752 656624
rect 86738 641952 98130 648996
rect 86738 641660 120688 641952
rect 136728 641660 148074 650176
rect 86738 641628 148074 641660
rect 151874 641628 353834 641660
rect 86738 641330 353834 641628
rect 402730 641404 404778 681322
rect 570592 646006 575942 683716
rect 565206 644560 576142 646006
rect 565206 641590 567706 644560
rect 431788 641404 433780 641410
rect 476622 641404 567706 641590
rect 86738 641284 362636 641330
rect 400454 641284 443936 641404
rect 86738 641242 443936 641284
rect 445822 641242 567706 641404
rect 86738 639756 567706 641242
rect 573760 639756 576142 644560
rect 86738 639526 576142 639756
rect 86738 633438 354208 639526
rect 360382 634562 576142 639526
rect 360382 633438 567668 634562
rect 86738 632060 567668 633438
rect 86738 631874 495080 632060
rect 86738 631718 362636 631874
rect 402730 631866 404778 631874
rect 86738 631234 353834 631718
rect 86738 631118 98130 631234
rect 116546 631184 353834 631234
rect 116546 631162 135504 631184
rect 151526 631162 353834 631184
rect 116546 631140 135360 631162
rect 186722 630690 191570 631162
rect 204138 630690 209704 631162
rect 186722 585092 191570 604984
rect 204138 591614 209704 604984
rect 204098 590968 209704 591614
rect 417434 592326 424178 631874
rect 565206 629758 567668 632060
rect 573722 629758 576142 634562
rect 565206 627532 576142 629758
rect 437706 592334 438460 592380
rect 437302 592326 438460 592334
rect 417434 592148 438460 592326
rect 417434 591984 437812 592148
rect 437996 591984 438212 592148
rect 438396 591984 438460 592148
rect 417434 591748 438460 591984
rect 417434 591584 437812 591748
rect 437996 591584 438212 591748
rect 438396 591584 438460 591748
rect 417434 591348 438460 591584
rect 417434 591184 437812 591348
rect 437996 591184 438212 591348
rect 438396 591184 438460 591348
rect 403550 591110 408774 591138
rect 403528 591104 408774 591110
rect 417434 591104 438460 591184
rect 204098 586508 209692 590968
rect 403528 590948 438460 591104
rect 403528 590784 437812 590948
rect 437996 590784 438212 590948
rect 438396 590784 438460 590948
rect 442320 592244 443082 592420
rect 446106 592378 446860 592380
rect 442320 592080 442412 592244
rect 442596 592080 442812 592244
rect 442996 592080 443082 592244
rect 442320 591918 443082 592080
rect 442320 591910 442760 591918
rect 442320 591606 442366 591910
rect 442650 591614 442760 591910
rect 443044 591614 443082 591918
rect 442650 591606 443082 591614
rect 442320 591444 443082 591606
rect 442320 591280 442412 591444
rect 442596 591280 442812 591444
rect 442996 591280 443082 591444
rect 442320 591126 443082 591280
rect 442320 590830 442356 591126
rect 442684 591122 443082 591126
rect 442684 590830 442768 591122
rect 442320 590818 442768 590830
rect 443052 590818 443082 591122
rect 442320 590816 443082 590818
rect 442324 590814 443082 590816
rect 445116 592148 446860 592378
rect 445116 591984 446212 592148
rect 446396 591984 446612 592148
rect 446796 591984 446860 592148
rect 445116 591748 446860 591984
rect 445116 591584 446212 591748
rect 446396 591584 446612 591748
rect 446796 591584 446860 591748
rect 445116 591348 446860 591584
rect 445116 591184 446212 591348
rect 446396 591184 446612 591348
rect 446796 591184 446860 591348
rect 445116 590948 446860 591184
rect 403528 590748 438460 590784
rect 403528 590732 437490 590748
rect 403528 590224 424178 590732
rect 403528 589642 424150 590224
rect 403528 588544 410472 589642
rect 411230 589624 424150 589642
rect 403528 588304 405560 588544
rect 405868 588304 406160 588544
rect 406468 588304 406760 588544
rect 407068 588304 407360 588544
rect 407668 588304 407960 588544
rect 408268 588304 408560 588544
rect 408868 588304 409160 588544
rect 409468 588304 410472 588544
rect 403528 588056 410472 588304
rect 417344 589300 424150 589624
rect 435922 589680 436970 590732
rect 437706 590720 438460 590748
rect 445116 590784 446212 590948
rect 446396 590784 446612 590948
rect 446796 590784 446860 590948
rect 450720 592244 451482 592420
rect 450720 592080 450812 592244
rect 450996 592080 451212 592244
rect 451396 592080 451482 592244
rect 450720 591918 451482 592080
rect 450720 591910 451160 591918
rect 450720 591606 450766 591910
rect 451050 591614 451160 591910
rect 451444 591614 451482 591918
rect 451050 591606 451482 591614
rect 450720 591444 451482 591606
rect 450720 591280 450812 591444
rect 450996 591280 451212 591444
rect 451396 591280 451482 591444
rect 450720 591126 451482 591280
rect 450720 590830 450756 591126
rect 451084 591122 451482 591126
rect 451084 590830 451168 591122
rect 450720 590818 451168 590830
rect 451452 590818 451482 591122
rect 450720 590816 451482 590818
rect 450724 590814 451482 590816
rect 445116 590720 446860 590784
rect 445116 589680 446108 590720
rect 417344 588084 424158 589300
rect 435922 588662 446108 589680
rect 403528 586456 404756 588056
rect 403528 586454 405494 586456
rect 403528 586344 410080 586454
rect 403528 586104 405560 586344
rect 405868 586104 406160 586344
rect 406468 586104 406760 586344
rect 407068 586104 407360 586344
rect 407668 586104 407960 586344
rect 408268 586104 408560 586344
rect 408868 586104 409160 586344
rect 409468 586104 410080 586344
rect 403528 586024 410080 586104
rect 416354 586336 417192 586444
rect 403528 586014 405494 586024
rect 416354 585948 416472 586336
rect 417092 585948 417192 586336
rect 416354 585850 417192 585948
rect 186716 584756 191570 585092
rect 416356 585216 417188 585316
rect 416356 584828 416474 585216
rect 417094 584828 417188 585216
rect 186716 584374 191564 584756
rect 416356 584730 417188 584828
rect 405234 581174 410146 581588
rect 405234 580628 405622 581174
rect 406400 580628 406822 581174
rect 407600 580628 408022 581174
rect 408800 580628 409222 581174
rect 410000 580628 410146 581174
rect 405234 580232 410146 580628
rect 141154 541976 150810 548702
<< via4 >>
rect 119008 695156 119292 695430
rect 67008 687156 67292 687430
rect 416166 687976 416450 688042
rect 416166 687812 416212 687976
rect 416212 687812 416396 687976
rect 416396 687812 416450 687976
rect 416166 687738 416450 687812
rect 416560 687976 416844 688050
rect 416560 687812 416612 687976
rect 416612 687812 416796 687976
rect 416796 687812 416844 687976
rect 416560 687746 416844 687812
rect 416156 687176 416484 687258
rect 416156 687012 416212 687176
rect 416212 687012 416396 687176
rect 416396 687012 416484 687176
rect 416156 686962 416484 687012
rect 416568 687176 416852 687254
rect 416568 687012 416622 687176
rect 416622 687012 416806 687176
rect 416806 687012 416852 687176
rect 416568 686950 416852 687012
rect 468166 687976 468450 688042
rect 468166 687812 468212 687976
rect 468212 687812 468396 687976
rect 468396 687812 468450 687976
rect 468166 687738 468450 687812
rect 468560 687976 468844 688050
rect 468560 687812 468612 687976
rect 468612 687812 468796 687976
rect 468796 687812 468844 687976
rect 468560 687746 468844 687812
rect 468156 687176 468484 687258
rect 468156 687012 468212 687176
rect 468212 687012 468396 687176
rect 468396 687012 468484 687176
rect 468156 686962 468484 687012
rect 468568 687176 468852 687254
rect 468568 687012 468622 687176
rect 468622 687012 468806 687176
rect 468806 687012 468852 687176
rect 468568 686950 468852 687012
rect 512924 686746 517294 691578
rect 519782 686746 524152 691578
rect 568166 687976 568450 688042
rect 568166 687812 568212 687976
rect 568212 687812 568396 687976
rect 568396 687812 568450 687976
rect 568166 687738 568450 687812
rect 568560 687976 568844 688050
rect 568560 687812 568612 687976
rect 568612 687812 568796 687976
rect 568796 687812 568844 687976
rect 568560 687746 568844 687812
rect 568156 687176 568484 687258
rect 568156 687012 568212 687176
rect 568212 687012 568396 687176
rect 568396 687012 568484 687176
rect 568156 686962 568484 687012
rect 568568 687176 568852 687254
rect 568568 687012 568622 687176
rect 568622 687012 568806 687176
rect 568806 687012 568852 687176
rect 568568 686950 568852 687012
rect 70008 673458 70292 673732
rect 121808 673220 122092 673494
rect 222764 656624 224356 664238
rect 442366 591844 442650 591910
rect 442366 591680 442412 591844
rect 442412 591680 442596 591844
rect 442596 591680 442650 591844
rect 442366 591606 442650 591680
rect 442760 591844 443044 591918
rect 442760 591680 442812 591844
rect 442812 591680 442996 591844
rect 442996 591680 443044 591844
rect 442760 591614 443044 591680
rect 442356 591044 442684 591126
rect 442356 590880 442412 591044
rect 442412 590880 442596 591044
rect 442596 590880 442684 591044
rect 442356 590830 442684 590880
rect 442768 591044 443052 591122
rect 442768 590880 442822 591044
rect 442822 590880 443006 591044
rect 443006 590880 443052 591044
rect 442768 590818 443052 590880
rect 450766 591844 451050 591910
rect 450766 591680 450812 591844
rect 450812 591680 450996 591844
rect 450996 591680 451050 591844
rect 450766 591606 451050 591680
rect 451160 591844 451444 591918
rect 451160 591680 451212 591844
rect 451212 591680 451396 591844
rect 451396 591680 451444 591844
rect 451160 591614 451444 591680
rect 450756 591044 451084 591126
rect 450756 590880 450812 591044
rect 450812 590880 450996 591044
rect 450996 590880 451084 591044
rect 450756 590830 451084 590880
rect 451168 591044 451452 591122
rect 451168 590880 451222 591044
rect 451222 590880 451406 591044
rect 451406 590880 451452 591044
rect 451168 590818 451452 590880
rect 416472 585948 417092 586336
rect 416474 584828 417094 585216
rect 405622 580628 406400 581174
rect 406822 580628 407600 581174
rect 408022 580628 408800 581174
rect 409222 580628 410000 581174
<< metal5 >>
rect 165594 700170 170596 704800
rect 175894 702300 180896 704800
rect 217294 702970 222294 704800
rect 217294 702300 222298 702970
rect 227594 702926 232594 704800
rect 175894 702254 180892 702300
rect 165578 698240 170596 700170
rect 44678 696132 54410 697566
rect 44678 695462 54460 696132
rect 44678 695454 116830 695462
rect 118970 695454 119334 695486
rect 44678 695430 119334 695454
rect 44678 695156 119008 695430
rect 119292 695156 119334 695430
rect 44678 695134 119334 695156
rect 44678 695062 116830 695134
rect 118970 695110 119334 695134
rect 44678 691616 54460 695062
rect 44804 687468 54460 691616
rect 44804 687454 66236 687468
rect 66970 687454 67334 687486
rect 44804 687430 67334 687454
rect 44804 687156 67008 687430
rect 67292 687156 67334 687430
rect 44804 687134 67334 687156
rect 44804 687126 66354 687134
rect 44804 687110 54468 687126
rect 66970 687110 67334 687134
rect 44804 673902 54460 687110
rect 165596 684280 170596 698240
rect 165600 682626 170596 684280
rect 175888 683670 180892 702254
rect 217306 700998 222298 702300
rect 217306 684124 222336 700998
rect 175908 682686 180892 683670
rect 175908 682660 187876 682686
rect 217280 682660 222336 684124
rect 227582 694624 232594 702926
rect 318994 702300 323994 704800
rect 329294 702300 334294 704800
rect 227582 682660 232548 694624
rect 511622 691578 524830 694392
rect 511622 689710 512924 691578
rect 416118 688050 416878 688698
rect 416118 688042 416560 688050
rect 416118 687738 416166 688042
rect 416450 687746 416560 688042
rect 416844 687850 416878 688050
rect 468118 688052 468878 688698
rect 473182 688052 474038 688056
rect 468118 688050 474038 688052
rect 468118 688042 468560 688050
rect 416844 687746 420894 687850
rect 416450 687738 420894 687746
rect 416118 687298 420894 687738
rect 416118 687258 416878 687298
rect 416118 686962 416156 687258
rect 416484 687254 416878 687258
rect 416484 686962 416568 687254
rect 416118 686950 416568 686962
rect 416852 686950 416878 687254
rect 416118 686838 416878 686950
rect 420072 686994 420894 687298
rect 468118 687738 468166 688042
rect 468450 687746 468560 688042
rect 468844 687746 474038 688050
rect 468450 687738 474038 687746
rect 468118 687500 474038 687738
rect 468118 687298 468896 687500
rect 468118 687258 468878 687298
rect 420072 685576 420916 686994
rect 468118 686962 468156 687258
rect 468484 687254 468878 687258
rect 468484 686962 468568 687254
rect 468118 686950 468568 686962
rect 468852 686950 468878 687254
rect 468118 686838 468878 686950
rect 473182 686592 474038 687500
rect 511498 686746 512924 689710
rect 517294 686746 519782 691578
rect 524152 689710 524830 691578
rect 566276 689710 568936 689756
rect 524152 688050 568936 689710
rect 524152 688042 568560 688050
rect 524152 687738 568166 688042
rect 568450 687746 568560 688042
rect 568844 687746 568936 688050
rect 568450 687738 568936 687746
rect 524152 687258 568936 687738
rect 524152 686962 568156 687258
rect 568484 687254 568936 687258
rect 568484 686962 568568 687254
rect 524152 686950 568568 686962
rect 568852 686950 568936 687254
rect 524152 686746 568936 686950
rect 175908 682658 191412 682660
rect 208250 682658 232548 682660
rect 175908 682626 191572 682658
rect 165600 677212 191572 682626
rect 175818 677200 181542 677212
rect 185920 677168 191572 677212
rect 44804 673888 66874 673902
rect 67330 673888 70382 673902
rect 44804 673732 70382 673888
rect 44804 673458 70008 673732
rect 70292 673458 70382 673732
rect 44804 673316 70382 673458
rect 44804 661200 54460 673316
rect 66380 673302 70382 673316
rect 103262 673632 111234 675078
rect 119710 673632 121470 673634
rect 103262 673494 122298 673632
rect 103262 673220 121808 673494
rect 122092 673220 122298 673494
rect 103262 673068 122298 673220
rect 44804 661186 99016 661200
rect 103262 661186 111234 673068
rect 44804 654946 111234 661186
rect 44804 653892 111288 654946
rect 44804 637908 54664 653892
rect 44908 630818 54664 637908
rect 44908 618130 54564 630818
rect 44908 613838 54488 618130
rect 44908 552254 54564 613838
rect 186724 585092 191572 677168
rect 204138 677168 232548 682658
rect 420086 681318 420914 685576
rect 265894 681262 420914 681318
rect 247820 681228 420914 681262
rect 473190 681228 474018 686592
rect 511498 686070 568936 686746
rect 511622 685510 568936 686070
rect 511622 681228 524830 685510
rect 566276 685486 568936 685510
rect 247820 677672 524916 681228
rect 247820 677366 524830 677672
rect 247820 677310 275360 677366
rect 419536 677340 524830 677366
rect 204138 591614 209704 677168
rect 222390 664238 224726 664668
rect 222390 656624 222764 664238
rect 224356 662136 224726 664238
rect 247820 662136 252154 677310
rect 224356 658694 252154 662136
rect 224356 656624 224726 658694
rect 247820 658682 252154 658694
rect 222390 656366 224726 656624
rect 443890 652480 445122 677340
rect 453350 652484 454564 677340
rect 443890 651668 445126 652480
rect 453350 652158 454576 652484
rect 443932 592430 445126 651668
rect 443228 592420 445126 592430
rect 453382 592426 454576 652158
rect 451650 592420 454582 592426
rect 204098 590968 209704 591614
rect 442316 591918 445126 592420
rect 442316 591910 442760 591918
rect 442316 591606 442366 591910
rect 442650 591614 442760 591910
rect 443044 591614 445126 591918
rect 442650 591606 445126 591614
rect 442316 591126 445126 591606
rect 204098 587862 209692 590968
rect 442316 590830 442356 591126
rect 442684 591122 445126 591126
rect 442684 590830 442768 591122
rect 442316 590818 442768 590830
rect 443052 590818 445126 591122
rect 442316 590732 445126 590818
rect 450716 591918 454582 592420
rect 450716 591910 451160 591918
rect 450716 591606 450766 591910
rect 451050 591614 451160 591910
rect 451444 591614 454582 591918
rect 451050 591606 454582 591614
rect 450716 591126 454582 591606
rect 450716 590830 450756 591126
rect 451084 591122 454582 591126
rect 451084 590830 451168 591122
rect 450716 590818 451168 590830
rect 451452 590818 454582 591122
rect 450716 590732 454582 590818
rect 443228 590724 445126 590732
rect 451650 590730 454582 590732
rect 443932 590722 445126 590724
rect 404884 587890 411558 587894
rect 416544 587890 416996 587892
rect 404360 587886 413436 587890
rect 415322 587886 416996 587890
rect 210580 587862 218504 587886
rect 230148 587862 416996 587886
rect 203986 587428 416996 587862
rect 203986 587396 417000 587428
rect 203986 587374 233540 587396
rect 404360 587384 413436 587396
rect 404884 587382 411780 587384
rect 404884 587380 411558 587382
rect 404894 587374 411558 587380
rect 416544 587374 417000 587396
rect 204098 586508 209692 587374
rect 416544 586444 417002 587374
rect 416354 586336 417192 586444
rect 416354 585948 416472 586336
rect 417092 585948 417192 586336
rect 416354 585850 417192 585948
rect 186718 584756 191572 585092
rect 416356 585216 417188 585316
rect 416356 584828 416474 585216
rect 417094 584828 417188 585216
rect 186718 583460 191566 584756
rect 416356 584730 417188 584828
rect 416576 583490 416994 584730
rect 409576 583468 416994 583490
rect 223086 583460 416994 583468
rect 186718 582996 416994 583460
rect 223086 582978 416994 582996
rect 409576 582974 416994 582978
rect 405234 581570 411694 581576
rect 417328 581570 425018 583368
rect 405234 581418 425018 581570
rect 405234 581174 424970 581418
rect 405234 580628 405622 581174
rect 406400 580628 406822 581174
rect 407600 580628 408022 581174
rect 408800 580628 409222 581174
rect 410000 580628 424970 581174
rect 405234 580238 424970 580628
rect 405234 580228 411694 580238
rect 417358 552254 424970 580238
rect 511622 554468 524830 677340
rect 44908 551998 434004 552254
rect 511624 552106 524830 554468
rect 44908 551888 476240 551998
rect 511624 551896 524886 552106
rect 499162 551888 524886 551896
rect 44908 542478 524886 551888
rect 44908 542110 434004 542478
rect 499162 542446 524886 542478
rect 44908 541976 54564 542110
<< comment >>
rect -100 704000 584100 704100
rect -100 0 0 704000
rect 584000 0 584100 704000
rect -100 -100 584100 0
use comparator_v6  comparator_v6_0
timestamp 1654337383
transform 0 1 419250 1 0 584722
box -2598 -1934 4390 5556
use sky130_fd_pr__diode_pd2nw_05v5_RT56W3  sky130_fd_pr__diode_pd2nw_05v5_RT56W3_0
timestamp 1654337383
transform 1 0 73460 0 1 687284
box -321 -321 321 321
use sky130_fd_pr__diode_pd2nw_05v5_RT56W3  sky130_fd_pr__diode_pd2nw_05v5_RT56W3_1
timestamp 1654337383
transform 1 0 125458 0 1 695284
box -321 -321 321 321
use sky130_fd_pr__diode_pw2nd_05v5_3P6M5Y  sky130_fd_pr__diode_pw2nd_05v5_3P6M5Y_0
timestamp 1654337383
transform 1 0 119582 0 1 695306
box -238 -238 238 238
use sky130_fd_pr__diode_pw2nd_05v5_GT7G3L  sky130_fd_pr__diode_pw2nd_05v5_GT7G3L_0
timestamp 1654337383
transform 1 0 67548 0 1 687302
box -183 -183 183 183
use sky130_fd_sc_hd__buf_2  sky130_fd_sc_hd__buf_2_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1654337383
transform 0 -1 440640 1 0 591294
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  sky130_fd_sc_hd__buf_2_1
timestamp 1654337383
transform 0 -1 448994 1 0 591314
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  sky130_fd_sc_hd__buf_2_2
timestamp 1654337383
transform 0 1 70516 -1 0 673768
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  sky130_fd_sc_hd__buf_2_3
timestamp 1654337383
transform 0 1 122500 -1 0 673516
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  sky130_fd_sc_hd__buf_2_4
timestamp 1654337383
transform 0 1 569338 -1 0 689064
box -38 -48 406 592
use sky130_fd_sc_hd__buf_16  sky130_fd_sc_hd__buf_16_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1654337383
transform 0 -1 415748 1 0 686664
box -38 -48 2062 592
use sky130_fd_sc_hd__buf_16  sky130_fd_sc_hd__buf_16_1
timestamp 1654337383
transform 0 -1 467556 1 0 686698
box -38 -48 2062 592
use sky130_fd_sc_hd__buf_16  sky130_fd_sc_hd__buf_16_2
timestamp 1654337383
transform 1 0 406656 0 1 587358
box -38 -48 2062 592
use sky130_fd_sc_hd__buf_16  sky130_fd_sc_hd__buf_16_3
timestamp 1654337383
transform 1 0 406646 0 1 585256
box -38 -48 2062 592
use sky130_fd_sc_hd__buf_16  sky130_fd_sc_hd__buf_16_4
timestamp 1654337383
transform 0 1 569338 -1 0 688388
box -38 -48 2062 592
<< labels >>
flabel metal3 s 582340 191430 584800 196230 0 FreeSans 1120 0 0 0 vssd1
port 568 nsew signal bidirectional
flabel metal3 s 582340 181430 584800 186230 0 FreeSans 1120 0 0 0 vssd1
port 569 nsew signal bidirectional
flabel metal2 s 6434 -800 6546 480 0 FreeSans 1120 90 0 0 wbs_we_i
port 677 nsew signal input
flabel metal2 s 5252 -800 5364 480 0 FreeSans 1120 90 0 0 wbs_stb_i
port 676 nsew signal input
flabel metal2 s 25346 -800 25458 480 0 FreeSans 1120 90 0 0 wbs_sel_i[3]
port 675 nsew signal input
flabel metal2 s 20618 -800 20730 480 0 FreeSans 1120 90 0 0 wbs_sel_i[2]
port 674 nsew signal input
flabel metal2 s 15890 -800 16002 480 0 FreeSans 1120 90 0 0 wbs_sel_i[1]
port 673 nsew signal input
flabel metal2 s 11162 -800 11274 480 0 FreeSans 1120 90 0 0 wbs_sel_i[0]
port 672 nsew signal input
flabel metal2 s 46622 -800 46734 480 0 FreeSans 1120 90 0 0 wbs_dat_o[9]
port 671 nsew signal tristate
flabel metal2 s 43076 -800 43188 480 0 FreeSans 1120 90 0 0 wbs_dat_o[8]
port 670 nsew signal tristate
flabel metal2 s 39530 -800 39642 480 0 FreeSans 1120 90 0 0 wbs_dat_o[7]
port 669 nsew signal tristate
flabel metal2 s 35984 -800 36096 480 0 FreeSans 1120 90 0 0 wbs_dat_o[6]
port 668 nsew signal tristate
flabel metal2 s 32438 -800 32550 480 0 FreeSans 1120 90 0 0 wbs_dat_o[5]
port 667 nsew signal tristate
flabel metal2 s 28892 -800 29004 480 0 FreeSans 1120 90 0 0 wbs_dat_o[4]
port 666 nsew signal tristate
flabel metal2 s 24164 -800 24276 480 0 FreeSans 1120 90 0 0 wbs_dat_o[3]
port 665 nsew signal tristate
flabel metal2 s 124634 -800 124746 480 0 FreeSans 1120 90 0 0 wbs_dat_o[31]
port 664 nsew signal tristate
flabel metal2 s 121088 -800 121200 480 0 FreeSans 1120 90 0 0 wbs_dat_o[30]
port 663 nsew signal tristate
flabel metal2 s 19436 -800 19548 480 0 FreeSans 1120 90 0 0 wbs_dat_o[2]
port 662 nsew signal tristate
flabel metal2 s 117542 -800 117654 480 0 FreeSans 1120 90 0 0 wbs_dat_o[29]
port 661 nsew signal tristate
flabel metal2 s 113996 -800 114108 480 0 FreeSans 1120 90 0 0 wbs_dat_o[28]
port 660 nsew signal tristate
flabel metal2 s 110450 -800 110562 480 0 FreeSans 1120 90 0 0 wbs_dat_o[27]
port 659 nsew signal tristate
flabel metal2 s 106904 -800 107016 480 0 FreeSans 1120 90 0 0 wbs_dat_o[26]
port 658 nsew signal tristate
flabel metal2 s 103358 -800 103470 480 0 FreeSans 1120 90 0 0 wbs_dat_o[25]
port 657 nsew signal tristate
flabel metal2 s 99812 -800 99924 480 0 FreeSans 1120 90 0 0 wbs_dat_o[24]
port 656 nsew signal tristate
flabel metal2 s 96266 -800 96378 480 0 FreeSans 1120 90 0 0 wbs_dat_o[23]
port 655 nsew signal tristate
flabel metal2 s 92720 -800 92832 480 0 FreeSans 1120 90 0 0 wbs_dat_o[22]
port 654 nsew signal tristate
flabel metal2 s 89174 -800 89286 480 0 FreeSans 1120 90 0 0 wbs_dat_o[21]
port 653 nsew signal tristate
flabel metal2 s 85628 -800 85740 480 0 FreeSans 1120 90 0 0 wbs_dat_o[20]
port 652 nsew signal tristate
flabel metal2 s 14708 -800 14820 480 0 FreeSans 1120 90 0 0 wbs_dat_o[1]
port 651 nsew signal tristate
flabel metal2 s 82082 -800 82194 480 0 FreeSans 1120 90 0 0 wbs_dat_o[19]
port 650 nsew signal tristate
flabel metal2 s 78536 -800 78648 480 0 FreeSans 1120 90 0 0 wbs_dat_o[18]
port 649 nsew signal tristate
flabel metal2 s 74990 -800 75102 480 0 FreeSans 1120 90 0 0 wbs_dat_o[17]
port 648 nsew signal tristate
flabel metal2 s 71444 -800 71556 480 0 FreeSans 1120 90 0 0 wbs_dat_o[16]
port 647 nsew signal tristate
flabel metal2 s 67898 -800 68010 480 0 FreeSans 1120 90 0 0 wbs_dat_o[15]
port 646 nsew signal tristate
flabel metal2 s 64352 -800 64464 480 0 FreeSans 1120 90 0 0 wbs_dat_o[14]
port 645 nsew signal tristate
flabel metal2 s 60806 -800 60918 480 0 FreeSans 1120 90 0 0 wbs_dat_o[13]
port 644 nsew signal tristate
flabel metal2 s 57260 -800 57372 480 0 FreeSans 1120 90 0 0 wbs_dat_o[12]
port 643 nsew signal tristate
flabel metal2 s 53714 -800 53826 480 0 FreeSans 1120 90 0 0 wbs_dat_o[11]
port 642 nsew signal tristate
flabel metal2 s 50168 -800 50280 480 0 FreeSans 1120 90 0 0 wbs_dat_o[10]
port 641 nsew signal tristate
flabel metal2 s 9980 -800 10092 480 0 FreeSans 1120 90 0 0 wbs_dat_o[0]
port 640 nsew signal tristate
flabel metal2 s 45440 -800 45552 480 0 FreeSans 1120 90 0 0 wbs_dat_i[9]
port 639 nsew signal input
flabel metal2 s 41894 -800 42006 480 0 FreeSans 1120 90 0 0 wbs_dat_i[8]
port 638 nsew signal input
flabel metal2 s 38348 -800 38460 480 0 FreeSans 1120 90 0 0 wbs_dat_i[7]
port 637 nsew signal input
flabel metal2 s 34802 -800 34914 480 0 FreeSans 1120 90 0 0 wbs_dat_i[6]
port 636 nsew signal input
flabel metal2 s 31256 -800 31368 480 0 FreeSans 1120 90 0 0 wbs_dat_i[5]
port 635 nsew signal input
flabel metal2 s 27710 -800 27822 480 0 FreeSans 1120 90 0 0 wbs_dat_i[4]
port 634 nsew signal input
flabel metal2 s 22982 -800 23094 480 0 FreeSans 1120 90 0 0 wbs_dat_i[3]
port 633 nsew signal input
flabel metal2 s 123452 -800 123564 480 0 FreeSans 1120 90 0 0 wbs_dat_i[31]
port 632 nsew signal input
flabel metal2 s 119906 -800 120018 480 0 FreeSans 1120 90 0 0 wbs_dat_i[30]
port 631 nsew signal input
flabel metal2 s 18254 -800 18366 480 0 FreeSans 1120 90 0 0 wbs_dat_i[2]
port 630 nsew signal input
flabel metal2 s 116360 -800 116472 480 0 FreeSans 1120 90 0 0 wbs_dat_i[29]
port 629 nsew signal input
flabel metal2 s 112814 -800 112926 480 0 FreeSans 1120 90 0 0 wbs_dat_i[28]
port 628 nsew signal input
flabel metal2 s 109268 -800 109380 480 0 FreeSans 1120 90 0 0 wbs_dat_i[27]
port 627 nsew signal input
flabel metal2 s 105722 -800 105834 480 0 FreeSans 1120 90 0 0 wbs_dat_i[26]
port 626 nsew signal input
flabel metal2 s 102176 -800 102288 480 0 FreeSans 1120 90 0 0 wbs_dat_i[25]
port 625 nsew signal input
flabel metal2 s 98630 -800 98742 480 0 FreeSans 1120 90 0 0 wbs_dat_i[24]
port 624 nsew signal input
flabel metal2 s 95084 -800 95196 480 0 FreeSans 1120 90 0 0 wbs_dat_i[23]
port 623 nsew signal input
flabel metal2 s 91538 -800 91650 480 0 FreeSans 1120 90 0 0 wbs_dat_i[22]
port 622 nsew signal input
flabel metal2 s 87992 -800 88104 480 0 FreeSans 1120 90 0 0 wbs_dat_i[21]
port 621 nsew signal input
flabel metal2 s 84446 -800 84558 480 0 FreeSans 1120 90 0 0 wbs_dat_i[20]
port 620 nsew signal input
flabel metal2 s 13526 -800 13638 480 0 FreeSans 1120 90 0 0 wbs_dat_i[1]
port 619 nsew signal input
flabel metal2 s 80900 -800 81012 480 0 FreeSans 1120 90 0 0 wbs_dat_i[19]
port 618 nsew signal input
flabel metal2 s 77354 -800 77466 480 0 FreeSans 1120 90 0 0 wbs_dat_i[18]
port 617 nsew signal input
flabel metal2 s 73808 -800 73920 480 0 FreeSans 1120 90 0 0 wbs_dat_i[17]
port 616 nsew signal input
flabel metal2 s 70262 -800 70374 480 0 FreeSans 1120 90 0 0 wbs_dat_i[16]
port 615 nsew signal input
flabel metal2 s 66716 -800 66828 480 0 FreeSans 1120 90 0 0 wbs_dat_i[15]
port 614 nsew signal input
flabel metal2 s 63170 -800 63282 480 0 FreeSans 1120 90 0 0 wbs_dat_i[14]
port 613 nsew signal input
flabel metal2 s 59624 -800 59736 480 0 FreeSans 1120 90 0 0 wbs_dat_i[13]
port 612 nsew signal input
flabel metal2 s 56078 -800 56190 480 0 FreeSans 1120 90 0 0 wbs_dat_i[12]
port 611 nsew signal input
flabel metal2 s 52532 -800 52644 480 0 FreeSans 1120 90 0 0 wbs_dat_i[11]
port 610 nsew signal input
flabel metal2 s 48986 -800 49098 480 0 FreeSans 1120 90 0 0 wbs_dat_i[10]
port 609 nsew signal input
flabel metal2 s 8798 -800 8910 480 0 FreeSans 1120 90 0 0 wbs_dat_i[0]
port 608 nsew signal input
flabel metal2 s 4070 -800 4182 480 0 FreeSans 1120 90 0 0 wbs_cyc_i
port 607 nsew signal input
flabel metal2 s 44258 -800 44370 480 0 FreeSans 1120 90 0 0 wbs_adr_i[9]
port 606 nsew signal input
flabel metal2 s 40712 -800 40824 480 0 FreeSans 1120 90 0 0 wbs_adr_i[8]
port 605 nsew signal input
flabel metal2 s 37166 -800 37278 480 0 FreeSans 1120 90 0 0 wbs_adr_i[7]
port 604 nsew signal input
flabel metal2 s 33620 -800 33732 480 0 FreeSans 1120 90 0 0 wbs_adr_i[6]
port 603 nsew signal input
flabel metal2 s 30074 -800 30186 480 0 FreeSans 1120 90 0 0 wbs_adr_i[5]
port 602 nsew signal input
flabel metal2 s 26528 -800 26640 480 0 FreeSans 1120 90 0 0 wbs_adr_i[4]
port 601 nsew signal input
flabel metal2 s 21800 -800 21912 480 0 FreeSans 1120 90 0 0 wbs_adr_i[3]
port 600 nsew signal input
flabel metal2 s 122270 -800 122382 480 0 FreeSans 1120 90 0 0 wbs_adr_i[31]
port 599 nsew signal input
flabel metal2 s 118724 -800 118836 480 0 FreeSans 1120 90 0 0 wbs_adr_i[30]
port 598 nsew signal input
flabel metal2 s 17072 -800 17184 480 0 FreeSans 1120 90 0 0 wbs_adr_i[2]
port 597 nsew signal input
flabel metal2 s 115178 -800 115290 480 0 FreeSans 1120 90 0 0 wbs_adr_i[29]
port 596 nsew signal input
flabel metal2 s 111632 -800 111744 480 0 FreeSans 1120 90 0 0 wbs_adr_i[28]
port 595 nsew signal input
flabel metal2 s 108086 -800 108198 480 0 FreeSans 1120 90 0 0 wbs_adr_i[27]
port 594 nsew signal input
flabel metal2 s 104540 -800 104652 480 0 FreeSans 1120 90 0 0 wbs_adr_i[26]
port 593 nsew signal input
flabel metal2 s 100994 -800 101106 480 0 FreeSans 1120 90 0 0 wbs_adr_i[25]
port 592 nsew signal input
flabel metal2 s 97448 -800 97560 480 0 FreeSans 1120 90 0 0 wbs_adr_i[24]
port 591 nsew signal input
flabel metal2 s 93902 -800 94014 480 0 FreeSans 1120 90 0 0 wbs_adr_i[23]
port 590 nsew signal input
flabel metal2 s 90356 -800 90468 480 0 FreeSans 1120 90 0 0 wbs_adr_i[22]
port 589 nsew signal input
flabel metal2 s 86810 -800 86922 480 0 FreeSans 1120 90 0 0 wbs_adr_i[21]
port 588 nsew signal input
flabel metal2 s 83264 -800 83376 480 0 FreeSans 1120 90 0 0 wbs_adr_i[20]
port 587 nsew signal input
flabel metal2 s 12344 -800 12456 480 0 FreeSans 1120 90 0 0 wbs_adr_i[1]
port 586 nsew signal input
flabel metal2 s 79718 -800 79830 480 0 FreeSans 1120 90 0 0 wbs_adr_i[19]
port 585 nsew signal input
flabel metal2 s 76172 -800 76284 480 0 FreeSans 1120 90 0 0 wbs_adr_i[18]
port 584 nsew signal input
flabel metal2 s 72626 -800 72738 480 0 FreeSans 1120 90 0 0 wbs_adr_i[17]
port 583 nsew signal input
flabel metal2 s 69080 -800 69192 480 0 FreeSans 1120 90 0 0 wbs_adr_i[16]
port 582 nsew signal input
flabel metal2 s 65534 -800 65646 480 0 FreeSans 1120 90 0 0 wbs_adr_i[15]
port 581 nsew signal input
flabel metal2 s 61988 -800 62100 480 0 FreeSans 1120 90 0 0 wbs_adr_i[14]
port 580 nsew signal input
flabel metal2 s 58442 -800 58554 480 0 FreeSans 1120 90 0 0 wbs_adr_i[13]
port 579 nsew signal input
flabel metal2 s 54896 -800 55008 480 0 FreeSans 1120 90 0 0 wbs_adr_i[12]
port 578 nsew signal input
flabel metal2 s 51350 -800 51462 480 0 FreeSans 1120 90 0 0 wbs_adr_i[11]
port 577 nsew signal input
flabel metal2 s 47804 -800 47916 480 0 FreeSans 1120 90 0 0 wbs_adr_i[10]
port 576 nsew signal input
flabel metal2 s 7616 -800 7728 480 0 FreeSans 1120 90 0 0 wbs_adr_i[0]
port 575 nsew signal input
flabel metal2 s 2888 -800 3000 480 0 FreeSans 1120 90 0 0 wbs_ack_o
port 574 nsew signal tristate
flabel metal2 s 1706 -800 1818 480 0 FreeSans 1120 90 0 0 wb_rst_i
port 573 nsew signal input
flabel metal2 s 524 -800 636 480 0 FreeSans 1120 90 0 0 wb_clk_i
port 572 nsew signal input
flabel metal3 s 0 162888 1660 167688 0 FreeSans 1120 0 0 0 vssd2
port 571 nsew signal bidirectional
flabel metal3 s 0 172888 1660 177688 0 FreeSans 1120 0 0 0 vssd2
port 570 nsew signal bidirectional
flabel metal3 s 0 549442 1660 554242 0 FreeSans 1120 0 0 0 vssa2
port 567 nsew signal bidirectional
flabel metal3 s 0 559442 1660 564242 0 FreeSans 1120 0 0 0 vssa2
port 566 nsew signal bidirectional
flabel metal3 s 582340 136830 584800 141630 0 FreeSans 1120 0 0 0 vssa1
port 565 nsew signal bidirectional
flabel metal3 s 582340 146830 584800 151630 0 FreeSans 1120 0 0 0 vssa1
port 564 nsew signal bidirectional
flabel metal3 s 510594 702340 515394 704800 0 FreeSans 1920 180 0 0 vssa1
port 563 nsew signal bidirectional
flabel metal3 s 520594 702340 525394 704800 0 FreeSans 1920 180 0 0 vssa1
port 562 nsew signal bidirectional
flabel metal3 s 0 214888 1660 219688 0 FreeSans 1120 0 0 0 vdda2
port 561 nsew signal bidirectional
flabel metal3 s 0 204888 1660 209688 0 FreeSans 1120 0 0 0 vdda2
port 560 nsew signal bidirectional
flabel metal3 s 582340 225230 584800 230030 0 FreeSans 1120 0 0 0 vdda1
port 559 nsew signal bidirectional
flabel metal3 s 582340 235230 584800 240030 0 FreeSans 1120 0 0 0 vdda1
port 558 nsew signal bidirectional
flabel metal3 s 582340 550562 584800 555362 0 FreeSans 1120 0 0 0 vdda1
port 557 nsew signal bidirectional
flabel metal3 s 582340 540562 584800 545362 0 FreeSans 1120 0 0 0 vdda1
port 556 nsew signal bidirectional
flabel metal3 s 0 633842 1660 638642 0 FreeSans 1120 0 0 0 vccd2
port 555 nsew signal bidirectional
flabel metal3 s 0 643842 1660 648642 0 FreeSans 1120 0 0 0 vccd2
port 554 nsew signal bidirectional
flabel metal3 s 582340 629784 584800 634584 0 FreeSans 1120 0 0 0 vccd1
port 553 nsew signal bidirectional
flabel metal3 s 582340 639784 584800 644584 0 FreeSans 1120 0 0 0 vccd1
port 552 nsew signal bidirectional
flabel metal2 s 583250 -800 583362 480 0 FreeSans 1120 90 0 0 user_irq[2]
port 551 nsew signal tristate
flabel metal2 s 582068 -800 582180 480 0 FreeSans 1120 90 0 0 user_irq[1]
port 550 nsew signal tristate
flabel metal2 s 580886 -800 580998 480 0 FreeSans 1120 90 0 0 user_irq[0]
port 549 nsew signal tristate
flabel metal2 s 579704 -800 579816 480 0 FreeSans 1120 90 0 0 user_clock2
port 548 nsew signal input
flabel metal2 s 160094 -800 160206 480 0 FreeSans 1120 90 0 0 la_oenb[9]
port 547 nsew signal input
flabel metal2 s 479234 -800 479346 480 0 FreeSans 1120 90 0 0 la_oenb[99]
port 546 nsew signal input
flabel metal2 s 475688 -800 475800 480 0 FreeSans 1120 90 0 0 la_oenb[98]
port 545 nsew signal input
flabel metal2 s 472142 -800 472254 480 0 FreeSans 1120 90 0 0 la_oenb[97]
port 544 nsew signal input
flabel metal2 s 468596 -800 468708 480 0 FreeSans 1120 90 0 0 la_oenb[96]
port 543 nsew signal input
flabel metal2 s 465050 -800 465162 480 0 FreeSans 1120 90 0 0 la_oenb[95]
port 542 nsew signal input
flabel metal2 s 461504 -800 461616 480 0 FreeSans 1120 90 0 0 la_oenb[94]
port 541 nsew signal input
flabel metal2 s 457958 -800 458070 480 0 FreeSans 1120 90 0 0 la_oenb[93]
port 540 nsew signal input
flabel metal2 s 454412 -800 454524 480 0 FreeSans 1120 90 0 0 la_oenb[92]
port 539 nsew signal input
flabel metal2 s 450866 -800 450978 480 0 FreeSans 1120 90 0 0 la_oenb[91]
port 538 nsew signal input
flabel metal2 s 447320 -800 447432 480 0 FreeSans 1120 90 0 0 la_oenb[90]
port 537 nsew signal input
flabel metal2 s 156548 -800 156660 480 0 FreeSans 1120 90 0 0 la_oenb[8]
port 536 nsew signal input
flabel metal2 s 443774 -800 443886 480 0 FreeSans 1120 90 0 0 la_oenb[89]
port 535 nsew signal input
flabel metal2 s 440228 -800 440340 480 0 FreeSans 1120 90 0 0 la_oenb[88]
port 534 nsew signal input
flabel metal2 s 436682 -800 436794 480 0 FreeSans 1120 90 0 0 la_oenb[87]
port 533 nsew signal input
flabel metal2 s 433136 -800 433248 480 0 FreeSans 1120 90 0 0 la_oenb[86]
port 532 nsew signal input
flabel metal2 s 429590 -800 429702 480 0 FreeSans 1120 90 0 0 la_oenb[85]
port 531 nsew signal input
flabel metal2 s 426044 -800 426156 480 0 FreeSans 1120 90 0 0 la_oenb[84]
port 530 nsew signal input
flabel metal2 s 422498 -800 422610 480 0 FreeSans 1120 90 0 0 la_oenb[83]
port 529 nsew signal input
flabel metal2 s 418952 -800 419064 480 0 FreeSans 1120 90 0 0 la_oenb[82]
port 528 nsew signal input
flabel metal2 s 415406 -800 415518 480 0 FreeSans 1120 90 0 0 la_oenb[81]
port 527 nsew signal input
flabel metal2 s 411860 -800 411972 480 0 FreeSans 1120 90 0 0 la_oenb[80]
port 526 nsew signal input
flabel metal2 s 153002 -800 153114 480 0 FreeSans 1120 90 0 0 la_oenb[7]
port 525 nsew signal input
flabel metal2 s 408314 -800 408426 480 0 FreeSans 1120 90 0 0 la_oenb[79]
port 524 nsew signal input
flabel metal2 s 404768 -800 404880 480 0 FreeSans 1120 90 0 0 la_oenb[78]
port 523 nsew signal input
flabel metal2 s 401222 -800 401334 480 0 FreeSans 1120 90 0 0 la_oenb[77]
port 522 nsew signal input
flabel metal2 s 397676 -800 397788 480 0 FreeSans 1120 90 0 0 la_oenb[76]
port 521 nsew signal input
flabel metal2 s 394130 -800 394242 480 0 FreeSans 1120 90 0 0 la_oenb[75]
port 520 nsew signal input
flabel metal2 s 390584 -800 390696 480 0 FreeSans 1120 90 0 0 la_oenb[74]
port 519 nsew signal input
flabel metal2 s 387038 -800 387150 480 0 FreeSans 1120 90 0 0 la_oenb[73]
port 518 nsew signal input
flabel metal2 s 383492 -800 383604 480 0 FreeSans 1120 90 0 0 la_oenb[72]
port 517 nsew signal input
flabel metal2 s 379946 -800 380058 480 0 FreeSans 1120 90 0 0 la_oenb[71]
port 516 nsew signal input
flabel metal2 s 376400 -800 376512 480 0 FreeSans 1120 90 0 0 la_oenb[70]
port 515 nsew signal input
flabel metal2 s 149456 -800 149568 480 0 FreeSans 1120 90 0 0 la_oenb[6]
port 514 nsew signal input
flabel metal2 s 372854 -800 372966 480 0 FreeSans 1120 90 0 0 la_oenb[69]
port 513 nsew signal input
flabel metal2 s 369308 -800 369420 480 0 FreeSans 1120 90 0 0 la_oenb[68]
port 512 nsew signal input
flabel metal2 s 365762 -800 365874 480 0 FreeSans 1120 90 0 0 la_oenb[67]
port 511 nsew signal input
flabel metal2 s 362216 -800 362328 480 0 FreeSans 1120 90 0 0 la_oenb[66]
port 510 nsew signal input
flabel metal2 s 358670 -800 358782 480 0 FreeSans 1120 90 0 0 la_oenb[65]
port 509 nsew signal input
flabel metal2 s 355124 -800 355236 480 0 FreeSans 1120 90 0 0 la_oenb[64]
port 508 nsew signal input
flabel metal2 s 351578 -800 351690 480 0 FreeSans 1120 90 0 0 la_oenb[63]
port 507 nsew signal input
flabel metal2 s 348032 -800 348144 480 0 FreeSans 1120 90 0 0 la_oenb[62]
port 506 nsew signal input
flabel metal2 s 344486 -800 344598 480 0 FreeSans 1120 90 0 0 la_oenb[61]
port 505 nsew signal input
flabel metal2 s 340940 -800 341052 480 0 FreeSans 1120 90 0 0 la_oenb[60]
port 504 nsew signal input
flabel metal2 s 145910 -800 146022 480 0 FreeSans 1120 90 0 0 la_oenb[5]
port 503 nsew signal input
flabel metal2 s 337394 -800 337506 480 0 FreeSans 1120 90 0 0 la_oenb[59]
port 502 nsew signal input
flabel metal2 s 333848 -800 333960 480 0 FreeSans 1120 90 0 0 la_oenb[58]
port 501 nsew signal input
flabel metal2 s 330302 -800 330414 480 0 FreeSans 1120 90 0 0 la_oenb[57]
port 500 nsew signal input
flabel metal2 s 326756 -800 326868 480 0 FreeSans 1120 90 0 0 la_oenb[56]
port 499 nsew signal input
flabel metal2 s 323210 -800 323322 480 0 FreeSans 1120 90 0 0 la_oenb[55]
port 498 nsew signal input
flabel metal2 s 319664 -800 319776 480 0 FreeSans 1120 90 0 0 la_oenb[54]
port 497 nsew signal input
flabel metal2 s 316118 -800 316230 480 0 FreeSans 1120 90 0 0 la_oenb[53]
port 496 nsew signal input
flabel metal2 s 312572 -800 312684 480 0 FreeSans 1120 90 0 0 la_oenb[52]
port 495 nsew signal input
flabel metal2 s 309026 -800 309138 480 0 FreeSans 1120 90 0 0 la_oenb[51]
port 494 nsew signal input
flabel metal2 s 305480 -800 305592 480 0 FreeSans 1120 90 0 0 la_oenb[50]
port 493 nsew signal input
flabel metal2 s 142364 -800 142476 480 0 FreeSans 1120 90 0 0 la_oenb[4]
port 492 nsew signal input
flabel metal2 s 301934 -800 302046 480 0 FreeSans 1120 90 0 0 la_oenb[49]
port 491 nsew signal input
flabel metal2 s 298388 -800 298500 480 0 FreeSans 1120 90 0 0 la_oenb[48]
port 490 nsew signal input
flabel metal2 s 294842 -800 294954 480 0 FreeSans 1120 90 0 0 la_oenb[47]
port 489 nsew signal input
flabel metal2 s 291296 -800 291408 480 0 FreeSans 1120 90 0 0 la_oenb[46]
port 488 nsew signal input
flabel metal2 s 287750 -800 287862 480 0 FreeSans 1120 90 0 0 la_oenb[45]
port 487 nsew signal input
flabel metal2 s 284204 -800 284316 480 0 FreeSans 1120 90 0 0 la_oenb[44]
port 486 nsew signal input
flabel metal2 s 280658 -800 280770 480 0 FreeSans 1120 90 0 0 la_oenb[43]
port 485 nsew signal input
flabel metal2 s 277112 -800 277224 480 0 FreeSans 1120 90 0 0 la_oenb[42]
port 484 nsew signal input
flabel metal2 s 273566 -800 273678 480 0 FreeSans 1120 90 0 0 la_oenb[41]
port 483 nsew signal input
flabel metal2 s 270020 -800 270132 480 0 FreeSans 1120 90 0 0 la_oenb[40]
port 482 nsew signal input
flabel metal2 s 138818 -800 138930 480 0 FreeSans 1120 90 0 0 la_oenb[3]
port 481 nsew signal input
flabel metal2 s 266474 -800 266586 480 0 FreeSans 1120 90 0 0 la_oenb[39]
port 480 nsew signal input
flabel metal2 s 262928 -800 263040 480 0 FreeSans 1120 90 0 0 la_oenb[38]
port 479 nsew signal input
flabel metal2 s 259382 -800 259494 480 0 FreeSans 1120 90 0 0 la_oenb[37]
port 478 nsew signal input
flabel metal2 s 255836 -800 255948 480 0 FreeSans 1120 90 0 0 la_oenb[36]
port 477 nsew signal input
flabel metal2 s 252290 -800 252402 480 0 FreeSans 1120 90 0 0 la_oenb[35]
port 476 nsew signal input
flabel metal2 s 248744 -800 248856 480 0 FreeSans 1120 90 0 0 la_oenb[34]
port 475 nsew signal input
flabel metal2 s 245198 -800 245310 480 0 FreeSans 1120 90 0 0 la_oenb[33]
port 474 nsew signal input
flabel metal2 s 241652 -800 241764 480 0 FreeSans 1120 90 0 0 la_oenb[32]
port 473 nsew signal input
flabel metal2 s 238106 -800 238218 480 0 FreeSans 1120 90 0 0 la_oenb[31]
port 472 nsew signal input
flabel metal2 s 234560 -800 234672 480 0 FreeSans 1120 90 0 0 la_oenb[30]
port 471 nsew signal input
flabel metal2 s 135272 -800 135384 480 0 FreeSans 1120 90 0 0 la_oenb[2]
port 470 nsew signal input
flabel metal2 s 231014 -800 231126 480 0 FreeSans 1120 90 0 0 la_oenb[29]
port 469 nsew signal input
flabel metal2 s 227468 -800 227580 480 0 FreeSans 1120 90 0 0 la_oenb[28]
port 468 nsew signal input
flabel metal2 s 223922 -800 224034 480 0 FreeSans 1120 90 0 0 la_oenb[27]
port 467 nsew signal input
flabel metal2 s 220376 -800 220488 480 0 FreeSans 1120 90 0 0 la_oenb[26]
port 466 nsew signal input
flabel metal2 s 216830 -800 216942 480 0 FreeSans 1120 90 0 0 la_oenb[25]
port 465 nsew signal input
flabel metal2 s 213284 -800 213396 480 0 FreeSans 1120 90 0 0 la_oenb[24]
port 464 nsew signal input
flabel metal2 s 209738 -800 209850 480 0 FreeSans 1120 90 0 0 la_oenb[23]
port 463 nsew signal input
flabel metal2 s 206192 -800 206304 480 0 FreeSans 1120 90 0 0 la_oenb[22]
port 462 nsew signal input
flabel metal2 s 202646 -800 202758 480 0 FreeSans 1120 90 0 0 la_oenb[21]
port 461 nsew signal input
flabel metal2 s 199100 -800 199212 480 0 FreeSans 1120 90 0 0 la_oenb[20]
port 460 nsew signal input
flabel metal2 s 131726 -800 131838 480 0 FreeSans 1120 90 0 0 la_oenb[1]
port 459 nsew signal input
flabel metal2 s 195554 -800 195666 480 0 FreeSans 1120 90 0 0 la_oenb[19]
port 458 nsew signal input
flabel metal2 s 192008 -800 192120 480 0 FreeSans 1120 90 0 0 la_oenb[18]
port 457 nsew signal input
flabel metal2 s 188462 -800 188574 480 0 FreeSans 1120 90 0 0 la_oenb[17]
port 456 nsew signal input
flabel metal2 s 184916 -800 185028 480 0 FreeSans 1120 90 0 0 la_oenb[16]
port 455 nsew signal input
flabel metal2 s 181370 -800 181482 480 0 FreeSans 1120 90 0 0 la_oenb[15]
port 454 nsew signal input
flabel metal2 s 177824 -800 177936 480 0 FreeSans 1120 90 0 0 la_oenb[14]
port 453 nsew signal input
flabel metal2 s 174278 -800 174390 480 0 FreeSans 1120 90 0 0 la_oenb[13]
port 452 nsew signal input
flabel metal2 s 170732 -800 170844 480 0 FreeSans 1120 90 0 0 la_oenb[12]
port 451 nsew signal input
flabel metal2 s 578522 -800 578634 480 0 FreeSans 1120 90 0 0 la_oenb[127]
port 450 nsew signal input
flabel metal2 s 574976 -800 575088 480 0 FreeSans 1120 90 0 0 la_oenb[126]
port 449 nsew signal input
flabel metal2 s 571430 -800 571542 480 0 FreeSans 1120 90 0 0 la_oenb[125]
port 448 nsew signal input
flabel metal2 s 567884 -800 567996 480 0 FreeSans 1120 90 0 0 la_oenb[124]
port 447 nsew signal input
flabel metal2 s 564338 -800 564450 480 0 FreeSans 1120 90 0 0 la_oenb[123]
port 446 nsew signal input
flabel metal2 s 560792 -800 560904 480 0 FreeSans 1120 90 0 0 la_oenb[122]
port 445 nsew signal input
flabel metal2 s 557246 -800 557358 480 0 FreeSans 1120 90 0 0 la_oenb[121]
port 444 nsew signal input
flabel metal2 s 553700 -800 553812 480 0 FreeSans 1120 90 0 0 la_oenb[120]
port 443 nsew signal input
flabel metal2 s 167186 -800 167298 480 0 FreeSans 1120 90 0 0 la_oenb[11]
port 442 nsew signal input
flabel metal2 s 550154 -800 550266 480 0 FreeSans 1120 90 0 0 la_oenb[119]
port 441 nsew signal input
flabel metal2 s 546608 -800 546720 480 0 FreeSans 1120 90 0 0 la_oenb[118]
port 440 nsew signal input
flabel metal2 s 543062 -800 543174 480 0 FreeSans 1120 90 0 0 la_oenb[117]
port 439 nsew signal input
flabel metal2 s 539516 -800 539628 480 0 FreeSans 1120 90 0 0 la_oenb[116]
port 438 nsew signal input
flabel metal2 s 535970 -800 536082 480 0 FreeSans 1120 90 0 0 la_oenb[115]
port 437 nsew signal input
flabel metal2 s 532424 -800 532536 480 0 FreeSans 1120 90 0 0 la_oenb[114]
port 436 nsew signal input
flabel metal2 s 528878 -800 528990 480 0 FreeSans 1120 90 0 0 la_oenb[113]
port 435 nsew signal input
flabel metal2 s 525332 -800 525444 480 0 FreeSans 1120 90 0 0 la_oenb[112]
port 434 nsew signal input
flabel metal2 s 521786 -800 521898 480 0 FreeSans 1120 90 0 0 la_oenb[111]
port 433 nsew signal input
flabel metal2 s 518240 -800 518352 480 0 FreeSans 1120 90 0 0 la_oenb[110]
port 432 nsew signal input
flabel metal2 s 163640 -800 163752 480 0 FreeSans 1120 90 0 0 la_oenb[10]
port 431 nsew signal input
flabel metal2 s 514694 -800 514806 480 0 FreeSans 1120 90 0 0 la_oenb[109]
port 430 nsew signal input
flabel metal2 s 511148 -800 511260 480 0 FreeSans 1120 90 0 0 la_oenb[108]
port 429 nsew signal input
flabel metal2 s 507602 -800 507714 480 0 FreeSans 1120 90 0 0 la_oenb[107]
port 428 nsew signal input
flabel metal2 s 504056 -800 504168 480 0 FreeSans 1120 90 0 0 la_oenb[106]
port 427 nsew signal input
flabel metal2 s 500510 -800 500622 480 0 FreeSans 1120 90 0 0 la_oenb[105]
port 426 nsew signal input
flabel metal2 s 496964 -800 497076 480 0 FreeSans 1120 90 0 0 la_oenb[104]
port 425 nsew signal input
flabel metal2 s 493418 -800 493530 480 0 FreeSans 1120 90 0 0 la_oenb[103]
port 424 nsew signal input
flabel metal2 s 489872 -800 489984 480 0 FreeSans 1120 90 0 0 la_oenb[102]
port 423 nsew signal input
flabel metal2 s 486326 -800 486438 480 0 FreeSans 1120 90 0 0 la_oenb[101]
port 422 nsew signal input
flabel metal2 s 482780 -800 482892 480 0 FreeSans 1120 90 0 0 la_oenb[100]
port 421 nsew signal input
flabel metal2 s 128180 -800 128292 480 0 FreeSans 1120 90 0 0 la_oenb[0]
port 420 nsew signal input
flabel metal2 s 158912 -800 159024 480 0 FreeSans 1120 90 0 0 la_data_out[9]
port 419 nsew signal tristate
flabel metal2 s 478052 -800 478164 480 0 FreeSans 1120 90 0 0 la_data_out[99]
port 418 nsew signal tristate
flabel metal2 s 474506 -800 474618 480 0 FreeSans 1120 90 0 0 la_data_out[98]
port 417 nsew signal tristate
flabel metal2 s 470960 -800 471072 480 0 FreeSans 1120 90 0 0 la_data_out[97]
port 416 nsew signal tristate
flabel metal2 s 467414 -800 467526 480 0 FreeSans 1120 90 0 0 la_data_out[96]
port 415 nsew signal tristate
flabel metal2 s 463868 -800 463980 480 0 FreeSans 1120 90 0 0 la_data_out[95]
port 414 nsew signal tristate
flabel metal2 s 460322 -800 460434 480 0 FreeSans 1120 90 0 0 la_data_out[94]
port 413 nsew signal tristate
flabel metal2 s 456776 -800 456888 480 0 FreeSans 1120 90 0 0 la_data_out[93]
port 412 nsew signal tristate
flabel metal2 s 453230 -800 453342 480 0 FreeSans 1120 90 0 0 la_data_out[92]
port 411 nsew signal tristate
flabel metal2 s 449684 -800 449796 480 0 FreeSans 1120 90 0 0 la_data_out[91]
port 410 nsew signal tristate
flabel metal2 s 446138 -800 446250 480 0 FreeSans 1120 90 0 0 la_data_out[90]
port 409 nsew signal tristate
flabel metal2 s 155366 -800 155478 480 0 FreeSans 1120 90 0 0 la_data_out[8]
port 408 nsew signal tristate
flabel metal2 s 442592 -800 442704 480 0 FreeSans 1120 90 0 0 la_data_out[89]
port 407 nsew signal tristate
flabel metal2 s 439046 -800 439158 480 0 FreeSans 1120 90 0 0 la_data_out[88]
port 406 nsew signal tristate
flabel metal2 s 435500 -800 435612 480 0 FreeSans 1120 90 0 0 la_data_out[87]
port 405 nsew signal tristate
flabel metal2 s 431954 -800 432066 480 0 FreeSans 1120 90 0 0 la_data_out[86]
port 404 nsew signal tristate
flabel metal2 s 428408 -800 428520 480 0 FreeSans 1120 90 0 0 la_data_out[85]
port 403 nsew signal tristate
flabel metal2 s 424862 -800 424974 480 0 FreeSans 1120 90 0 0 la_data_out[84]
port 402 nsew signal tristate
flabel metal2 s 421316 -800 421428 480 0 FreeSans 1120 90 0 0 la_data_out[83]
port 401 nsew signal tristate
flabel metal2 s 417770 -800 417882 480 0 FreeSans 1120 90 0 0 la_data_out[82]
port 400 nsew signal tristate
flabel metal2 s 414224 -800 414336 480 0 FreeSans 1120 90 0 0 la_data_out[81]
port 399 nsew signal tristate
flabel metal2 s 410678 -800 410790 480 0 FreeSans 1120 90 0 0 la_data_out[80]
port 398 nsew signal tristate
flabel metal2 s 151820 -800 151932 480 0 FreeSans 1120 90 0 0 la_data_out[7]
port 397 nsew signal tristate
flabel metal2 s 407132 -800 407244 480 0 FreeSans 1120 90 0 0 la_data_out[79]
port 396 nsew signal tristate
flabel metal2 s 403586 -800 403698 480 0 FreeSans 1120 90 0 0 la_data_out[78]
port 395 nsew signal tristate
flabel metal2 s 400040 -800 400152 480 0 FreeSans 1120 90 0 0 la_data_out[77]
port 394 nsew signal tristate
flabel metal2 s 396494 -800 396606 480 0 FreeSans 1120 90 0 0 la_data_out[76]
port 393 nsew signal tristate
flabel metal2 s 392948 -800 393060 480 0 FreeSans 1120 90 0 0 la_data_out[75]
port 392 nsew signal tristate
flabel metal2 s 389402 -800 389514 480 0 FreeSans 1120 90 0 0 la_data_out[74]
port 391 nsew signal tristate
flabel metal2 s 385856 -800 385968 480 0 FreeSans 1120 90 0 0 la_data_out[73]
port 390 nsew signal tristate
flabel metal2 s 382310 -800 382422 480 0 FreeSans 1120 90 0 0 la_data_out[72]
port 389 nsew signal tristate
flabel metal2 s 378764 -800 378876 480 0 FreeSans 1120 90 0 0 la_data_out[71]
port 388 nsew signal tristate
flabel metal2 s 375218 -800 375330 480 0 FreeSans 1120 90 0 0 la_data_out[70]
port 387 nsew signal tristate
flabel metal2 s 148274 -800 148386 480 0 FreeSans 1120 90 0 0 la_data_out[6]
port 386 nsew signal tristate
flabel metal2 s 371672 -800 371784 480 0 FreeSans 1120 90 0 0 la_data_out[69]
port 385 nsew signal tristate
flabel metal2 s 368126 -800 368238 480 0 FreeSans 1120 90 0 0 la_data_out[68]
port 384 nsew signal tristate
flabel metal2 s 364580 -800 364692 480 0 FreeSans 1120 90 0 0 la_data_out[67]
port 383 nsew signal tristate
flabel metal2 s 361034 -800 361146 480 0 FreeSans 1120 90 0 0 la_data_out[66]
port 382 nsew signal tristate
flabel metal2 s 357488 -800 357600 480 0 FreeSans 1120 90 0 0 la_data_out[65]
port 381 nsew signal tristate
flabel metal2 s 353942 -800 354054 480 0 FreeSans 1120 90 0 0 la_data_out[64]
port 380 nsew signal tristate
flabel metal2 s 350396 -800 350508 480 0 FreeSans 1120 90 0 0 la_data_out[63]
port 379 nsew signal tristate
flabel metal2 s 346850 -800 346962 480 0 FreeSans 1120 90 0 0 la_data_out[62]
port 378 nsew signal tristate
flabel metal2 s 343304 -800 343416 480 0 FreeSans 1120 90 0 0 la_data_out[61]
port 377 nsew signal tristate
flabel metal2 s 339758 -800 339870 480 0 FreeSans 1120 90 0 0 la_data_out[60]
port 376 nsew signal tristate
flabel metal2 s 144728 -800 144840 480 0 FreeSans 1120 90 0 0 la_data_out[5]
port 375 nsew signal tristate
flabel metal2 s 336212 -800 336324 480 0 FreeSans 1120 90 0 0 la_data_out[59]
port 374 nsew signal tristate
flabel metal2 s 332666 -800 332778 480 0 FreeSans 1120 90 0 0 la_data_out[58]
port 373 nsew signal tristate
flabel metal2 s 329120 -800 329232 480 0 FreeSans 1120 90 0 0 la_data_out[57]
port 372 nsew signal tristate
flabel metal2 s 325574 -800 325686 480 0 FreeSans 1120 90 0 0 la_data_out[56]
port 371 nsew signal tristate
flabel metal2 s 322028 -800 322140 480 0 FreeSans 1120 90 0 0 la_data_out[55]
port 370 nsew signal tristate
flabel metal2 s 318482 -800 318594 480 0 FreeSans 1120 90 0 0 la_data_out[54]
port 369 nsew signal tristate
flabel metal2 s 314936 -800 315048 480 0 FreeSans 1120 90 0 0 la_data_out[53]
port 368 nsew signal tristate
flabel metal2 s 311390 -800 311502 480 0 FreeSans 1120 90 0 0 la_data_out[52]
port 367 nsew signal tristate
flabel metal2 s 307844 -800 307956 480 0 FreeSans 1120 90 0 0 la_data_out[51]
port 366 nsew signal tristate
flabel metal2 s 304298 -800 304410 480 0 FreeSans 1120 90 0 0 la_data_out[50]
port 365 nsew signal tristate
flabel metal2 s 141182 -800 141294 480 0 FreeSans 1120 90 0 0 la_data_out[4]
port 364 nsew signal tristate
flabel metal2 s 300752 -800 300864 480 0 FreeSans 1120 90 0 0 la_data_out[49]
port 363 nsew signal tristate
flabel metal2 s 297206 -800 297318 480 0 FreeSans 1120 90 0 0 la_data_out[48]
port 362 nsew signal tristate
flabel metal2 s 293660 -800 293772 480 0 FreeSans 1120 90 0 0 la_data_out[47]
port 361 nsew signal tristate
flabel metal2 s 290114 -800 290226 480 0 FreeSans 1120 90 0 0 la_data_out[46]
port 360 nsew signal tristate
flabel metal2 s 286568 -800 286680 480 0 FreeSans 1120 90 0 0 la_data_out[45]
port 359 nsew signal tristate
flabel metal2 s 283022 -800 283134 480 0 FreeSans 1120 90 0 0 la_data_out[44]
port 358 nsew signal tristate
flabel metal2 s 279476 -800 279588 480 0 FreeSans 1120 90 0 0 la_data_out[43]
port 357 nsew signal tristate
flabel metal2 s 275930 -800 276042 480 0 FreeSans 1120 90 0 0 la_data_out[42]
port 356 nsew signal tristate
flabel metal2 s 272384 -800 272496 480 0 FreeSans 1120 90 0 0 la_data_out[41]
port 355 nsew signal tristate
flabel metal2 s 268838 -800 268950 480 0 FreeSans 1120 90 0 0 la_data_out[40]
port 354 nsew signal tristate
flabel metal2 s 137636 -800 137748 480 0 FreeSans 1120 90 0 0 la_data_out[3]
port 353 nsew signal tristate
flabel metal2 s 265292 -800 265404 480 0 FreeSans 1120 90 0 0 la_data_out[39]
port 352 nsew signal tristate
flabel metal2 s 261746 -800 261858 480 0 FreeSans 1120 90 0 0 la_data_out[38]
port 351 nsew signal tristate
flabel metal2 s 258200 -800 258312 480 0 FreeSans 1120 90 0 0 la_data_out[37]
port 350 nsew signal tristate
flabel metal2 s 254654 -800 254766 480 0 FreeSans 1120 90 0 0 la_data_out[36]
port 349 nsew signal tristate
flabel metal2 s 251108 -800 251220 480 0 FreeSans 1120 90 0 0 la_data_out[35]
port 348 nsew signal tristate
flabel metal2 s 247562 -800 247674 480 0 FreeSans 1120 90 0 0 la_data_out[34]
port 347 nsew signal tristate
flabel metal2 s 244016 -800 244128 480 0 FreeSans 1120 90 0 0 la_data_out[33]
port 346 nsew signal tristate
flabel metal2 s 240470 -800 240582 480 0 FreeSans 1120 90 0 0 la_data_out[32]
port 345 nsew signal tristate
flabel metal2 s 236924 -800 237036 480 0 FreeSans 1120 90 0 0 la_data_out[31]
port 344 nsew signal tristate
flabel metal2 s 233378 -800 233490 480 0 FreeSans 1120 90 0 0 la_data_out[30]
port 343 nsew signal tristate
flabel metal2 s 134090 -800 134202 480 0 FreeSans 1120 90 0 0 la_data_out[2]
port 342 nsew signal tristate
flabel metal2 s 229832 -800 229944 480 0 FreeSans 1120 90 0 0 la_data_out[29]
port 341 nsew signal tristate
flabel metal2 s 226286 -800 226398 480 0 FreeSans 1120 90 0 0 la_data_out[28]
port 340 nsew signal tristate
flabel metal2 s 222740 -800 222852 480 0 FreeSans 1120 90 0 0 la_data_out[27]
port 339 nsew signal tristate
flabel metal2 s 219194 -800 219306 480 0 FreeSans 1120 90 0 0 la_data_out[26]
port 338 nsew signal tristate
flabel metal2 s 215648 -800 215760 480 0 FreeSans 1120 90 0 0 la_data_out[25]
port 337 nsew signal tristate
flabel metal2 s 212102 -800 212214 480 0 FreeSans 1120 90 0 0 la_data_out[24]
port 336 nsew signal tristate
flabel metal2 s 208556 -800 208668 480 0 FreeSans 1120 90 0 0 la_data_out[23]
port 335 nsew signal tristate
flabel metal2 s 205010 -800 205122 480 0 FreeSans 1120 90 0 0 la_data_out[22]
port 334 nsew signal tristate
flabel metal2 s 201464 -800 201576 480 0 FreeSans 1120 90 0 0 la_data_out[21]
port 333 nsew signal tristate
flabel metal2 s 197918 -800 198030 480 0 FreeSans 1120 90 0 0 la_data_out[20]
port 332 nsew signal tristate
flabel metal2 s 130544 -800 130656 480 0 FreeSans 1120 90 0 0 la_data_out[1]
port 331 nsew signal tristate
flabel metal2 s 194372 -800 194484 480 0 FreeSans 1120 90 0 0 la_data_out[19]
port 330 nsew signal tristate
flabel metal2 s 190826 -800 190938 480 0 FreeSans 1120 90 0 0 la_data_out[18]
port 329 nsew signal tristate
flabel metal2 s 187280 -800 187392 480 0 FreeSans 1120 90 0 0 la_data_out[17]
port 328 nsew signal tristate
flabel metal2 s 183734 -800 183846 480 0 FreeSans 1120 90 0 0 la_data_out[16]
port 327 nsew signal tristate
flabel metal2 s 180188 -800 180300 480 0 FreeSans 1120 90 0 0 la_data_out[15]
port 326 nsew signal tristate
flabel metal2 s 176642 -800 176754 480 0 FreeSans 1120 90 0 0 la_data_out[14]
port 325 nsew signal tristate
flabel metal2 s 173096 -800 173208 480 0 FreeSans 1120 90 0 0 la_data_out[13]
port 324 nsew signal tristate
flabel metal2 s 169550 -800 169662 480 0 FreeSans 1120 90 0 0 la_data_out[12]
port 323 nsew signal tristate
flabel metal2 s 577340 -800 577452 480 0 FreeSans 1120 90 0 0 la_data_out[127]
port 322 nsew signal tristate
flabel metal2 s 573794 -800 573906 480 0 FreeSans 1120 90 0 0 la_data_out[126]
port 321 nsew signal tristate
flabel metal2 s 570248 -800 570360 480 0 FreeSans 1120 90 0 0 la_data_out[125]
port 320 nsew signal tristate
flabel metal2 s 566702 -800 566814 480 0 FreeSans 1120 90 0 0 la_data_out[124]
port 319 nsew signal tristate
flabel metal2 s 563156 -800 563268 480 0 FreeSans 1120 90 0 0 la_data_out[123]
port 318 nsew signal tristate
flabel metal2 s 559610 -800 559722 480 0 FreeSans 1120 90 0 0 la_data_out[122]
port 317 nsew signal tristate
flabel metal2 s 556064 -800 556176 480 0 FreeSans 1120 90 0 0 la_data_out[121]
port 316 nsew signal tristate
flabel metal2 s 552518 -800 552630 480 0 FreeSans 1120 90 0 0 la_data_out[120]
port 315 nsew signal tristate
flabel metal2 s 166004 -800 166116 480 0 FreeSans 1120 90 0 0 la_data_out[11]
port 314 nsew signal tristate
flabel metal2 s 548972 -800 549084 480 0 FreeSans 1120 90 0 0 la_data_out[119]
port 313 nsew signal tristate
flabel metal2 s 545426 -800 545538 480 0 FreeSans 1120 90 0 0 la_data_out[118]
port 312 nsew signal tristate
flabel metal2 s 541880 -800 541992 480 0 FreeSans 1120 90 0 0 la_data_out[117]
port 311 nsew signal tristate
flabel metal2 s 538334 -800 538446 480 0 FreeSans 1120 90 0 0 la_data_out[116]
port 310 nsew signal tristate
flabel metal2 s 534788 -800 534900 480 0 FreeSans 1120 90 0 0 la_data_out[115]
port 309 nsew signal tristate
flabel metal2 s 531242 -800 531354 480 0 FreeSans 1120 90 0 0 la_data_out[114]
port 308 nsew signal tristate
flabel metal2 s 527696 -800 527808 480 0 FreeSans 1120 90 0 0 la_data_out[113]
port 307 nsew signal tristate
flabel metal2 s 524150 -800 524262 480 0 FreeSans 1120 90 0 0 la_data_out[112]
port 306 nsew signal tristate
flabel metal2 s 520604 -800 520716 480 0 FreeSans 1120 90 0 0 la_data_out[111]
port 305 nsew signal tristate
flabel metal2 s 517058 -800 517170 480 0 FreeSans 1120 90 0 0 la_data_out[110]
port 304 nsew signal tristate
flabel metal2 s 162458 -800 162570 480 0 FreeSans 1120 90 0 0 la_data_out[10]
port 303 nsew signal tristate
flabel metal2 s 513512 -800 513624 480 0 FreeSans 1120 90 0 0 la_data_out[109]
port 302 nsew signal tristate
flabel metal2 s 509966 -800 510078 480 0 FreeSans 1120 90 0 0 la_data_out[108]
port 301 nsew signal tristate
flabel metal2 s 506420 -800 506532 480 0 FreeSans 1120 90 0 0 la_data_out[107]
port 300 nsew signal tristate
flabel metal2 s 502874 -800 502986 480 0 FreeSans 1120 90 0 0 la_data_out[106]
port 299 nsew signal tristate
flabel metal2 s 499328 -800 499440 480 0 FreeSans 1120 90 0 0 la_data_out[105]
port 298 nsew signal tristate
flabel metal2 s 495782 -800 495894 480 0 FreeSans 1120 90 0 0 la_data_out[104]
port 297 nsew signal tristate
flabel metal2 s 492236 -800 492348 480 0 FreeSans 1120 90 0 0 la_data_out[103]
port 296 nsew signal tristate
flabel metal2 s 488690 -800 488802 480 0 FreeSans 1120 90 0 0 la_data_out[102]
port 295 nsew signal tristate
flabel metal2 s 485144 -800 485256 480 0 FreeSans 1120 90 0 0 la_data_out[101]
port 294 nsew signal tristate
flabel metal2 s 481598 -800 481710 480 0 FreeSans 1120 90 0 0 la_data_out[100]
port 293 nsew signal tristate
flabel metal2 s 126998 -800 127110 480 0 FreeSans 1120 90 0 0 la_data_out[0]
port 292 nsew signal tristate
flabel metal2 s 157730 -800 157842 480 0 FreeSans 1120 90 0 0 la_data_in[9]
port 291 nsew signal input
flabel metal2 s 476870 -800 476982 480 0 FreeSans 1120 90 0 0 la_data_in[99]
port 290 nsew signal input
flabel metal2 s 473324 -800 473436 480 0 FreeSans 1120 90 0 0 la_data_in[98]
port 289 nsew signal input
flabel metal2 s 469778 -800 469890 480 0 FreeSans 1120 90 0 0 la_data_in[97]
port 288 nsew signal input
flabel metal2 s 466232 -800 466344 480 0 FreeSans 1120 90 0 0 la_data_in[96]
port 287 nsew signal input
flabel metal2 s 462686 -800 462798 480 0 FreeSans 1120 90 0 0 la_data_in[95]
port 286 nsew signal input
flabel metal2 s 459140 -800 459252 480 0 FreeSans 1120 90 0 0 la_data_in[94]
port 285 nsew signal input
flabel metal2 s 455594 -800 455706 480 0 FreeSans 1120 90 0 0 la_data_in[93]
port 284 nsew signal input
flabel metal2 s 452048 -800 452160 480 0 FreeSans 1120 90 0 0 la_data_in[92]
port 283 nsew signal input
flabel metal2 s 448502 -800 448614 480 0 FreeSans 1120 90 0 0 la_data_in[91]
port 282 nsew signal input
flabel metal2 s 444956 -800 445068 480 0 FreeSans 1120 90 0 0 la_data_in[90]
port 281 nsew signal input
flabel metal2 s 154184 -800 154296 480 0 FreeSans 1120 90 0 0 la_data_in[8]
port 280 nsew signal input
flabel metal2 s 441410 -800 441522 480 0 FreeSans 1120 90 0 0 la_data_in[89]
port 279 nsew signal input
flabel metal2 s 437864 -800 437976 480 0 FreeSans 1120 90 0 0 la_data_in[88]
port 278 nsew signal input
flabel metal2 s 434318 -800 434430 480 0 FreeSans 1120 90 0 0 la_data_in[87]
port 277 nsew signal input
flabel metal2 s 430772 -800 430884 480 0 FreeSans 1120 90 0 0 la_data_in[86]
port 276 nsew signal input
flabel metal2 s 427226 -800 427338 480 0 FreeSans 1120 90 0 0 la_data_in[85]
port 275 nsew signal input
flabel metal2 s 423680 -800 423792 480 0 FreeSans 1120 90 0 0 la_data_in[84]
port 274 nsew signal input
flabel metal2 s 420134 -800 420246 480 0 FreeSans 1120 90 0 0 la_data_in[83]
port 273 nsew signal input
flabel metal2 s 416588 -800 416700 480 0 FreeSans 1120 90 0 0 la_data_in[82]
port 272 nsew signal input
flabel metal2 s 413042 -800 413154 480 0 FreeSans 1120 90 0 0 la_data_in[81]
port 271 nsew signal input
flabel metal2 s 409496 -800 409608 480 0 FreeSans 1120 90 0 0 la_data_in[80]
port 270 nsew signal input
flabel metal2 s 150638 -800 150750 480 0 FreeSans 1120 90 0 0 la_data_in[7]
port 269 nsew signal input
flabel metal2 s 405950 -800 406062 480 0 FreeSans 1120 90 0 0 la_data_in[79]
port 268 nsew signal input
flabel metal2 s 402404 -800 402516 480 0 FreeSans 1120 90 0 0 la_data_in[78]
port 267 nsew signal input
flabel metal2 s 398858 -800 398970 480 0 FreeSans 1120 90 0 0 la_data_in[77]
port 266 nsew signal input
flabel metal2 s 395312 -800 395424 480 0 FreeSans 1120 90 0 0 la_data_in[76]
port 265 nsew signal input
flabel metal2 s 391766 -800 391878 480 0 FreeSans 1120 90 0 0 la_data_in[75]
port 264 nsew signal input
flabel metal2 s 388220 -800 388332 480 0 FreeSans 1120 90 0 0 la_data_in[74]
port 263 nsew signal input
flabel metal2 s 384674 -800 384786 480 0 FreeSans 1120 90 0 0 la_data_in[73]
port 262 nsew signal input
flabel metal2 s 381128 -800 381240 480 0 FreeSans 1120 90 0 0 la_data_in[72]
port 261 nsew signal input
flabel metal2 s 377582 -800 377694 480 0 FreeSans 1120 90 0 0 la_data_in[71]
port 260 nsew signal input
flabel metal2 s 374036 -800 374148 480 0 FreeSans 1120 90 0 0 la_data_in[70]
port 259 nsew signal input
flabel metal2 s 147092 -800 147204 480 0 FreeSans 1120 90 0 0 la_data_in[6]
port 258 nsew signal input
flabel metal2 s 370490 -800 370602 480 0 FreeSans 1120 90 0 0 la_data_in[69]
port 257 nsew signal input
flabel metal2 s 366944 -800 367056 480 0 FreeSans 1120 90 0 0 la_data_in[68]
port 256 nsew signal input
flabel metal2 s 363398 -800 363510 480 0 FreeSans 1120 90 0 0 la_data_in[67]
port 255 nsew signal input
flabel metal2 s 359852 -800 359964 480 0 FreeSans 1120 90 0 0 la_data_in[66]
port 254 nsew signal input
flabel metal2 s 356306 -800 356418 480 0 FreeSans 1120 90 0 0 la_data_in[65]
port 253 nsew signal input
flabel metal2 s 352760 -800 352872 480 0 FreeSans 1120 90 0 0 la_data_in[64]
port 252 nsew signal input
flabel metal2 s 349214 -800 349326 480 0 FreeSans 1120 90 0 0 la_data_in[63]
port 251 nsew signal input
flabel metal2 s 345668 -800 345780 480 0 FreeSans 1120 90 0 0 la_data_in[62]
port 250 nsew signal input
flabel metal2 s 342122 -800 342234 480 0 FreeSans 1120 90 0 0 la_data_in[61]
port 249 nsew signal input
flabel metal2 s 338576 -800 338688 480 0 FreeSans 1120 90 0 0 la_data_in[60]
port 248 nsew signal input
flabel metal2 s 143546 -800 143658 480 0 FreeSans 1120 90 0 0 la_data_in[5]
port 247 nsew signal input
flabel metal2 s 335030 -800 335142 480 0 FreeSans 1120 90 0 0 la_data_in[59]
port 246 nsew signal input
flabel metal2 s 331484 -800 331596 480 0 FreeSans 1120 90 0 0 la_data_in[58]
port 245 nsew signal input
flabel metal2 s 327938 -800 328050 480 0 FreeSans 1120 90 0 0 la_data_in[57]
port 244 nsew signal input
flabel metal2 s 324392 -800 324504 480 0 FreeSans 1120 90 0 0 la_data_in[56]
port 243 nsew signal input
flabel metal2 s 320846 -800 320958 480 0 FreeSans 1120 90 0 0 la_data_in[55]
port 242 nsew signal input
flabel metal2 s 317300 -800 317412 480 0 FreeSans 1120 90 0 0 la_data_in[54]
port 241 nsew signal input
flabel metal2 s 313754 -800 313866 480 0 FreeSans 1120 90 0 0 la_data_in[53]
port 240 nsew signal input
flabel metal2 s 310208 -800 310320 480 0 FreeSans 1120 90 0 0 la_data_in[52]
port 239 nsew signal input
flabel metal2 s 306662 -800 306774 480 0 FreeSans 1120 90 0 0 la_data_in[51]
port 238 nsew signal input
flabel metal2 s 303116 -800 303228 480 0 FreeSans 1120 90 0 0 la_data_in[50]
port 237 nsew signal input
flabel metal2 s 140000 -800 140112 480 0 FreeSans 1120 90 0 0 la_data_in[4]
port 236 nsew signal input
flabel metal2 s 299570 -800 299682 480 0 FreeSans 1120 90 0 0 la_data_in[49]
port 235 nsew signal input
flabel metal2 s 296024 -800 296136 480 0 FreeSans 1120 90 0 0 la_data_in[48]
port 234 nsew signal input
flabel metal2 s 292478 -800 292590 480 0 FreeSans 1120 90 0 0 la_data_in[47]
port 233 nsew signal input
flabel metal2 s 288932 -800 289044 480 0 FreeSans 1120 90 0 0 la_data_in[46]
port 232 nsew signal input
flabel metal2 s 285386 -800 285498 480 0 FreeSans 1120 90 0 0 la_data_in[45]
port 231 nsew signal input
flabel metal2 s 281840 -800 281952 480 0 FreeSans 1120 90 0 0 la_data_in[44]
port 230 nsew signal input
flabel metal2 s 278294 -800 278406 480 0 FreeSans 1120 90 0 0 la_data_in[43]
port 229 nsew signal input
flabel metal2 s 274748 -800 274860 480 0 FreeSans 1120 90 0 0 la_data_in[42]
port 228 nsew signal input
flabel metal2 s 271202 -800 271314 480 0 FreeSans 1120 90 0 0 la_data_in[41]
port 227 nsew signal input
flabel metal2 s 267656 -800 267768 480 0 FreeSans 1120 90 0 0 la_data_in[40]
port 226 nsew signal input
flabel metal2 s 136454 -800 136566 480 0 FreeSans 1120 90 0 0 la_data_in[3]
port 225 nsew signal input
flabel metal2 s 264110 -800 264222 480 0 FreeSans 1120 90 0 0 la_data_in[39]
port 224 nsew signal input
flabel metal2 s 260564 -800 260676 480 0 FreeSans 1120 90 0 0 la_data_in[38]
port 223 nsew signal input
flabel metal2 s 257018 -800 257130 480 0 FreeSans 1120 90 0 0 la_data_in[37]
port 222 nsew signal input
flabel metal2 s 253472 -800 253584 480 0 FreeSans 1120 90 0 0 la_data_in[36]
port 221 nsew signal input
flabel metal2 s 249926 -800 250038 480 0 FreeSans 1120 90 0 0 la_data_in[35]
port 220 nsew signal input
flabel metal2 s 246380 -800 246492 480 0 FreeSans 1120 90 0 0 la_data_in[34]
port 219 nsew signal input
flabel metal2 s 242834 -800 242946 480 0 FreeSans 1120 90 0 0 la_data_in[33]
port 218 nsew signal input
flabel metal2 s 239288 -800 239400 480 0 FreeSans 1120 90 0 0 la_data_in[32]
port 217 nsew signal input
flabel metal2 s 235742 -800 235854 480 0 FreeSans 1120 90 0 0 la_data_in[31]
port 216 nsew signal input
flabel metal2 s 232196 -800 232308 480 0 FreeSans 1120 90 0 0 la_data_in[30]
port 215 nsew signal input
flabel metal2 s 132908 -800 133020 480 0 FreeSans 1120 90 0 0 la_data_in[2]
port 214 nsew signal input
flabel metal2 s 228650 -800 228762 480 0 FreeSans 1120 90 0 0 la_data_in[29]
port 213 nsew signal input
flabel metal2 s 225104 -800 225216 480 0 FreeSans 1120 90 0 0 la_data_in[28]
port 212 nsew signal input
flabel metal2 s 221558 -800 221670 480 0 FreeSans 1120 90 0 0 la_data_in[27]
port 211 nsew signal input
flabel metal2 s 218012 -800 218124 480 0 FreeSans 1120 90 0 0 la_data_in[26]
port 210 nsew signal input
flabel metal2 s 214466 -800 214578 480 0 FreeSans 1120 90 0 0 la_data_in[25]
port 209 nsew signal input
flabel metal2 s 210920 -800 211032 480 0 FreeSans 1120 90 0 0 la_data_in[24]
port 208 nsew signal input
flabel metal2 s 207374 -800 207486 480 0 FreeSans 1120 90 0 0 la_data_in[23]
port 207 nsew signal input
flabel metal2 s 203828 -800 203940 480 0 FreeSans 1120 90 0 0 la_data_in[22]
port 206 nsew signal input
flabel metal2 s 200282 -800 200394 480 0 FreeSans 1120 90 0 0 la_data_in[21]
port 205 nsew signal input
flabel metal2 s 196736 -800 196848 480 0 FreeSans 1120 90 0 0 la_data_in[20]
port 204 nsew signal input
flabel metal2 s 129362 -800 129474 480 0 FreeSans 1120 90 0 0 la_data_in[1]
port 203 nsew signal input
flabel metal2 s 193190 -800 193302 480 0 FreeSans 1120 90 0 0 la_data_in[19]
port 202 nsew signal input
flabel metal2 s 189644 -800 189756 480 0 FreeSans 1120 90 0 0 la_data_in[18]
port 201 nsew signal input
flabel metal2 s 186098 -800 186210 480 0 FreeSans 1120 90 0 0 la_data_in[17]
port 200 nsew signal input
flabel metal2 s 182552 -800 182664 480 0 FreeSans 1120 90 0 0 la_data_in[16]
port 199 nsew signal input
flabel metal2 s 179006 -800 179118 480 0 FreeSans 1120 90 0 0 la_data_in[15]
port 198 nsew signal input
flabel metal2 s 175460 -800 175572 480 0 FreeSans 1120 90 0 0 la_data_in[14]
port 197 nsew signal input
flabel metal2 s 171914 -800 172026 480 0 FreeSans 1120 90 0 0 la_data_in[13]
port 196 nsew signal input
flabel metal2 s 168368 -800 168480 480 0 FreeSans 1120 90 0 0 la_data_in[12]
port 195 nsew signal input
flabel metal2 s 576158 -800 576270 480 0 FreeSans 1120 90 0 0 la_data_in[127]
port 194 nsew signal input
flabel metal2 s 572612 -800 572724 480 0 FreeSans 1120 90 0 0 la_data_in[126]
port 193 nsew signal input
flabel metal2 s 569066 -800 569178 480 0 FreeSans 1120 90 0 0 la_data_in[125]
port 192 nsew signal input
flabel metal2 s 565520 -800 565632 480 0 FreeSans 1120 90 0 0 la_data_in[124]
port 191 nsew signal input
flabel metal2 s 561974 -800 562086 480 0 FreeSans 1120 90 0 0 la_data_in[123]
port 190 nsew signal input
flabel metal2 s 558428 -800 558540 480 0 FreeSans 1120 90 0 0 la_data_in[122]
port 189 nsew signal input
flabel metal2 s 554882 -800 554994 480 0 FreeSans 1120 90 0 0 la_data_in[121]
port 188 nsew signal input
flabel metal2 s 551336 -800 551448 480 0 FreeSans 1120 90 0 0 la_data_in[120]
port 187 nsew signal input
flabel metal2 s 164822 -800 164934 480 0 FreeSans 1120 90 0 0 la_data_in[11]
port 186 nsew signal input
flabel metal2 s 547790 -800 547902 480 0 FreeSans 1120 90 0 0 la_data_in[119]
port 185 nsew signal input
flabel metal2 s 544244 -800 544356 480 0 FreeSans 1120 90 0 0 la_data_in[118]
port 184 nsew signal input
flabel metal2 s 540698 -800 540810 480 0 FreeSans 1120 90 0 0 la_data_in[117]
port 183 nsew signal input
flabel metal2 s 537152 -800 537264 480 0 FreeSans 1120 90 0 0 la_data_in[116]
port 182 nsew signal input
flabel metal2 s 533606 -800 533718 480 0 FreeSans 1120 90 0 0 la_data_in[115]
port 181 nsew signal input
flabel metal2 s 530060 -800 530172 480 0 FreeSans 1120 90 0 0 la_data_in[114]
port 180 nsew signal input
flabel metal2 s 526514 -800 526626 480 0 FreeSans 1120 90 0 0 la_data_in[113]
port 179 nsew signal input
flabel metal2 s 522968 -800 523080 480 0 FreeSans 1120 90 0 0 la_data_in[112]
port 178 nsew signal input
flabel metal2 s 519422 -800 519534 480 0 FreeSans 1120 90 0 0 la_data_in[111]
port 177 nsew signal input
flabel metal2 s 515876 -800 515988 480 0 FreeSans 1120 90 0 0 la_data_in[110]
port 176 nsew signal input
flabel metal2 s 161276 -800 161388 480 0 FreeSans 1120 90 0 0 la_data_in[10]
port 175 nsew signal input
flabel metal2 s 512330 -800 512442 480 0 FreeSans 1120 90 0 0 la_data_in[109]
port 174 nsew signal input
flabel metal2 s 508784 -800 508896 480 0 FreeSans 1120 90 0 0 la_data_in[108]
port 173 nsew signal input
flabel metal2 s 505238 -800 505350 480 0 FreeSans 1120 90 0 0 la_data_in[107]
port 172 nsew signal input
flabel metal2 s 501692 -800 501804 480 0 FreeSans 1120 90 0 0 la_data_in[106]
port 171 nsew signal input
flabel metal2 s 498146 -800 498258 480 0 FreeSans 1120 90 0 0 la_data_in[105]
port 170 nsew signal input
flabel metal2 s 494600 -800 494712 480 0 FreeSans 1120 90 0 0 la_data_in[104]
port 169 nsew signal input
flabel metal2 s 491054 -800 491166 480 0 FreeSans 1120 90 0 0 la_data_in[103]
port 168 nsew signal input
flabel metal2 s 487508 -800 487620 480 0 FreeSans 1120 90 0 0 la_data_in[102]
port 167 nsew signal input
flabel metal2 s 483962 -800 484074 480 0 FreeSans 1120 90 0 0 la_data_in[101]
port 166 nsew signal input
flabel metal2 s 480416 -800 480528 480 0 FreeSans 1120 90 0 0 la_data_in[100]
port 165 nsew signal input
flabel metal2 s 125816 -800 125928 480 0 FreeSans 1120 90 0 0 la_data_in[0]
port 164 nsew signal input
flabel metal3 s 583520 363602 584800 363714 0 FreeSans 1120 0 0 0 io_out[9]
port 163 nsew signal tristate
flabel metal3 s 583520 318380 584800 318492 0 FreeSans 1120 0 0 0 io_out[8]
port 162 nsew signal tristate
flabel metal3 s 583520 273958 584800 274070 0 FreeSans 1120 0 0 0 io_out[7]
port 161 nsew signal tristate
flabel metal3 s 583520 93936 584800 94048 0 FreeSans 1120 0 0 0 io_out[6]
port 160 nsew signal tristate
flabel metal3 s 583520 49278 584800 49390 0 FreeSans 1120 0 0 0 io_out[5]
port 159 nsew signal tristate
flabel metal3 s 583520 22820 584800 22932 0 FreeSans 1120 0 0 0 io_out[4]
port 158 nsew signal tristate
flabel metal3 s 583520 18092 584800 18204 0 FreeSans 1120 0 0 0 io_out[3]
port 157 nsew signal tristate
flabel metal3 s 583520 13364 584800 13476 0 FreeSans 1120 0 0 0 io_out[2]
port 156 nsew signal tristate
flabel metal3 s -800 2726 480 2838 0 FreeSans 1120 0 0 0 io_out[26]
port 155 nsew signal tristate
flabel metal3 s -800 7454 480 7566 0 FreeSans 1120 0 0 0 io_out[25]
port 154 nsew signal tristate
flabel metal3 s -800 12182 480 12294 0 FreeSans 1120 0 0 0 io_out[24]
port 153 nsew signal tristate
flabel metal3 s -800 33604 480 33716 0 FreeSans 1120 0 0 0 io_out[23]
port 152 nsew signal tristate
flabel metal3 s -800 76826 480 76938 0 FreeSans 1120 0 0 0 io_out[22]
port 151 nsew signal tristate
flabel metal3 s -800 120048 480 120160 0 FreeSans 1120 0 0 0 io_out[21]
port 150 nsew signal tristate
flabel metal3 s -800 247670 480 247782 0 FreeSans 1120 0 0 0 io_out[20]
port 149 nsew signal tristate
flabel metal3 s 583520 8636 584800 8748 0 FreeSans 1120 0 0 0 io_out[1]
port 148 nsew signal tristate
flabel metal3 s -800 290692 480 290804 0 FreeSans 1120 0 0 0 io_out[19]
port 147 nsew signal tristate
flabel metal3 s -800 333914 480 334026 0 FreeSans 1120 0 0 0 io_out[18]
port 146 nsew signal tristate
flabel metal3 s -800 377136 480 377248 0 FreeSans 1120 0 0 0 io_out[17]
port 145 nsew signal tristate
flabel metal3 s -800 420358 480 420470 0 FreeSans 1120 0 0 0 io_out[16]
port 144 nsew signal tristate
flabel metal3 s -800 463580 480 463692 0 FreeSans 1120 0 0 0 io_out[15]
port 143 nsew signal tristate
flabel metal3 s -800 506802 480 506914 0 FreeSans 1120 0 0 0 io_out[14]
port 142 nsew signal tristate
flabel metal3 s 583520 588290 584800 588402 0 FreeSans 1120 0 0 0 io_out[13]
port 141 nsew signal tristate
flabel metal3 s 583520 498868 584800 498980 0 FreeSans 1120 0 0 0 io_out[12]
port 140 nsew signal tristate
flabel metal3 s 583520 454446 584800 454558 0 FreeSans 1120 0 0 0 io_out[11]
port 139 nsew signal tristate
flabel metal3 s 583520 410024 584800 410136 0 FreeSans 1120 0 0 0 io_out[10]
port 138 nsew signal tristate
flabel metal3 s 583520 3908 584800 4020 0 FreeSans 1120 0 0 0 io_out[0]
port 137 nsew signal tristate
flabel metal3 s 583520 364784 584800 364896 0 FreeSans 1120 0 0 0 io_oeb[9]
port 136 nsew signal tristate
flabel metal3 s 583520 319562 584800 319674 0 FreeSans 1120 0 0 0 io_oeb[8]
port 135 nsew signal tristate
flabel metal3 s 583520 275140 584800 275252 0 FreeSans 1120 0 0 0 io_oeb[7]
port 134 nsew signal tristate
flabel metal3 s 583520 95118 584800 95230 0 FreeSans 1120 0 0 0 io_oeb[6]
port 133 nsew signal tristate
flabel metal3 s 583520 50460 584800 50572 0 FreeSans 1120 0 0 0 io_oeb[5]
port 132 nsew signal tristate
flabel metal3 s 583520 24002 584800 24114 0 FreeSans 1120 0 0 0 io_oeb[4]
port 131 nsew signal tristate
flabel metal3 s 583520 19274 584800 19386 0 FreeSans 1120 0 0 0 io_oeb[3]
port 130 nsew signal tristate
flabel metal3 s 583520 14546 584800 14658 0 FreeSans 1120 0 0 0 io_oeb[2]
port 129 nsew signal tristate
flabel metal3 s -800 1544 480 1656 0 FreeSans 1120 0 0 0 io_oeb[26]
port 128 nsew signal tristate
flabel metal3 s -800 6272 480 6384 0 FreeSans 1120 0 0 0 io_oeb[25]
port 127 nsew signal tristate
flabel metal3 s -800 11000 480 11112 0 FreeSans 1120 0 0 0 io_oeb[24]
port 126 nsew signal tristate
flabel metal3 s -800 32422 480 32534 0 FreeSans 1120 0 0 0 io_oeb[23]
port 125 nsew signal tristate
flabel metal3 s -800 75644 480 75756 0 FreeSans 1120 0 0 0 io_oeb[22]
port 124 nsew signal tristate
flabel metal3 s -800 118866 480 118978 0 FreeSans 1120 0 0 0 io_oeb[21]
port 123 nsew signal tristate
flabel metal3 s -800 246488 480 246600 0 FreeSans 1120 0 0 0 io_oeb[20]
port 122 nsew signal tristate
flabel metal3 s 583520 9818 584800 9930 0 FreeSans 1120 0 0 0 io_oeb[1]
port 121 nsew signal tristate
flabel metal3 s -800 289510 480 289622 0 FreeSans 1120 0 0 0 io_oeb[19]
port 120 nsew signal tristate
flabel metal3 s -800 332732 480 332844 0 FreeSans 1120 0 0 0 io_oeb[18]
port 119 nsew signal tristate
flabel metal3 s -800 375954 480 376066 0 FreeSans 1120 0 0 0 io_oeb[17]
port 118 nsew signal tristate
flabel metal3 s -800 419176 480 419288 0 FreeSans 1120 0 0 0 io_oeb[16]
port 117 nsew signal tristate
flabel metal3 s -800 462398 480 462510 0 FreeSans 1120 0 0 0 io_oeb[15]
port 116 nsew signal tristate
flabel metal3 s -800 505620 480 505732 0 FreeSans 1120 0 0 0 io_oeb[14]
port 115 nsew signal tristate
flabel metal3 s 583520 589472 584800 589584 0 FreeSans 1120 0 0 0 io_oeb[13]
port 114 nsew signal tristate
flabel metal3 s 583520 500050 584800 500162 0 FreeSans 1120 0 0 0 io_oeb[12]
port 113 nsew signal tristate
flabel metal3 s 583520 455628 584800 455740 0 FreeSans 1120 0 0 0 io_oeb[11]
port 112 nsew signal tristate
flabel metal3 s 583520 411206 584800 411318 0 FreeSans 1120 0 0 0 io_oeb[10]
port 111 nsew signal tristate
flabel metal3 s 583520 5090 584800 5202 0 FreeSans 1120 0 0 0 io_oeb[0]
port 110 nsew signal tristate
flabel metal3 s 583520 361238 584800 361350 0 FreeSans 1120 0 0 0 io_in_3v3[9]
port 109 nsew signal input
flabel metal3 s 583520 316016 584800 316128 0 FreeSans 1120 0 0 0 io_in_3v3[8]
port 108 nsew signal input
flabel metal3 s 583520 271594 584800 271706 0 FreeSans 1120 0 0 0 io_in_3v3[7]
port 107 nsew signal input
flabel metal3 s 583520 91572 584800 91684 0 FreeSans 1120 0 0 0 io_in_3v3[6]
port 106 nsew signal input
flabel metal3 s 583520 46914 584800 47026 0 FreeSans 1120 0 0 0 io_in_3v3[5]
port 105 nsew signal input
flabel metal3 s 583520 20456 584800 20568 0 FreeSans 1120 0 0 0 io_in_3v3[4]
port 104 nsew signal input
flabel metal3 s 583520 15728 584800 15840 0 FreeSans 1120 0 0 0 io_in_3v3[3]
port 103 nsew signal input
flabel metal3 s 583520 11000 584800 11112 0 FreeSans 1120 0 0 0 io_in_3v3[2]
port 102 nsew signal input
flabel metal3 s -800 5090 480 5202 0 FreeSans 1120 0 0 0 io_in_3v3[26]
port 101 nsew signal input
flabel metal3 s -800 9818 480 9930 0 FreeSans 1120 0 0 0 io_in_3v3[25]
port 100 nsew signal input
flabel metal3 s -800 14546 480 14658 0 FreeSans 1120 0 0 0 io_in_3v3[24]
port 99 nsew signal input
flabel metal3 s -800 35968 480 36080 0 FreeSans 1120 0 0 0 io_in_3v3[23]
port 98 nsew signal input
flabel metal3 s -800 79190 480 79302 0 FreeSans 1120 0 0 0 io_in_3v3[22]
port 97 nsew signal input
flabel metal3 s -800 122412 480 122524 0 FreeSans 1120 0 0 0 io_in_3v3[21]
port 96 nsew signal input
flabel metal3 s -800 250034 480 250146 0 FreeSans 1120 0 0 0 io_in_3v3[20]
port 95 nsew signal input
flabel metal3 s 583520 6272 584800 6384 0 FreeSans 1120 0 0 0 io_in_3v3[1]
port 94 nsew signal input
flabel metal3 s -800 293056 480 293168 0 FreeSans 1120 0 0 0 io_in_3v3[19]
port 93 nsew signal input
flabel metal3 s -800 336278 480 336390 0 FreeSans 1120 0 0 0 io_in_3v3[18]
port 92 nsew signal input
flabel metal3 s -800 379500 480 379612 0 FreeSans 1120 0 0 0 io_in_3v3[17]
port 91 nsew signal input
flabel metal3 s -800 422722 480 422834 0 FreeSans 1120 0 0 0 io_in_3v3[16]
port 90 nsew signal input
flabel metal3 s -800 465944 480 466056 0 FreeSans 1120 0 0 0 io_in_3v3[15]
port 89 nsew signal input
flabel metal3 s -800 509166 480 509278 0 FreeSans 1120 0 0 0 io_in_3v3[14]
port 88 nsew signal input
flabel metal3 s 583520 585926 584800 586038 0 FreeSans 1120 0 0 0 io_in_3v3[13]
port 87 nsew signal input
flabel metal3 s 583520 496504 584800 496616 0 FreeSans 1120 0 0 0 io_in_3v3[12]
port 86 nsew signal input
flabel metal3 s 583520 452082 584800 452194 0 FreeSans 1120 0 0 0 io_in_3v3[11]
port 85 nsew signal input
flabel metal3 s 583520 407660 584800 407772 0 FreeSans 1120 0 0 0 io_in_3v3[10]
port 84 nsew signal input
flabel metal3 s 583520 1544 584800 1656 0 FreeSans 1120 0 0 0 io_in_3v3[0]
port 83 nsew signal input
flabel metal3 s 583520 362420 584800 362532 0 FreeSans 1120 0 0 0 io_in[9]
port 82 nsew signal input
flabel metal3 s 583520 317198 584800 317310 0 FreeSans 1120 0 0 0 io_in[8]
port 81 nsew signal input
flabel metal3 s 583520 272776 584800 272888 0 FreeSans 1120 0 0 0 io_in[7]
port 80 nsew signal input
flabel metal3 s 583520 92754 584800 92866 0 FreeSans 1120 0 0 0 io_in[6]
port 79 nsew signal input
flabel metal3 s 583520 48096 584800 48208 0 FreeSans 1120 0 0 0 io_in[5]
port 78 nsew signal input
flabel metal3 s 583520 21638 584800 21750 0 FreeSans 1120 0 0 0 io_in[4]
port 77 nsew signal input
flabel metal3 s 583520 16910 584800 17022 0 FreeSans 1120 0 0 0 io_in[3]
port 76 nsew signal input
flabel metal3 s 583520 12182 584800 12294 0 FreeSans 1120 0 0 0 io_in[2]
port 75 nsew signal input
flabel metal3 s -800 3908 480 4020 0 FreeSans 1120 0 0 0 io_in[26]
port 74 nsew signal input
flabel metal3 s -800 8636 480 8748 0 FreeSans 1120 0 0 0 io_in[25]
port 73 nsew signal input
flabel metal3 s -800 13364 480 13476 0 FreeSans 1120 0 0 0 io_in[24]
port 72 nsew signal input
flabel metal3 s -800 34786 480 34898 0 FreeSans 1120 0 0 0 io_in[23]
port 71 nsew signal input
flabel metal3 s -800 78008 480 78120 0 FreeSans 1120 0 0 0 io_in[22]
port 70 nsew signal input
flabel metal3 s -800 121230 480 121342 0 FreeSans 1120 0 0 0 io_in[21]
port 69 nsew signal input
flabel metal3 s -800 248852 480 248964 0 FreeSans 1120 0 0 0 io_in[20]
port 68 nsew signal input
flabel metal3 s 583520 7454 584800 7566 0 FreeSans 1120 0 0 0 io_in[1]
port 67 nsew signal input
flabel metal3 s -800 291874 480 291986 0 FreeSans 1120 0 0 0 io_in[19]
port 66 nsew signal input
flabel metal3 s -800 335096 480 335208 0 FreeSans 1120 0 0 0 io_in[18]
port 65 nsew signal input
flabel metal3 s -800 378318 480 378430 0 FreeSans 1120 0 0 0 io_in[17]
port 64 nsew signal input
flabel metal3 s -800 421540 480 421652 0 FreeSans 1120 0 0 0 io_in[16]
port 63 nsew signal input
flabel metal3 s -800 464762 480 464874 0 FreeSans 1120 0 0 0 io_in[15]
port 62 nsew signal input
flabel metal3 s -800 507984 480 508096 0 FreeSans 1120 0 0 0 io_in[14]
port 61 nsew signal input
flabel metal3 s 583520 587108 584800 587220 0 FreeSans 1120 0 0 0 io_in[13]
port 60 nsew signal input
flabel metal3 s 583520 497686 584800 497798 0 FreeSans 1120 0 0 0 io_in[12]
port 59 nsew signal input
flabel metal3 s 583520 453264 584800 453376 0 FreeSans 1120 0 0 0 io_in[11]
port 58 nsew signal input
flabel metal3 s 583520 408842 584800 408954 0 FreeSans 1120 0 0 0 io_in[10]
port 57 nsew signal input
flabel metal3 s 583520 2726 584800 2838 0 FreeSans 1120 0 0 0 io_in[0]
port 56 nsew signal input
flabel metal3 s 170894 702300 173094 704800 0 FreeSans 1920 180 0 0 io_clamp_low[2]
port 55 nsew signal bidirectional
flabel metal3 s 222594 702300 224794 704800 0 FreeSans 1920 180 0 0 io_clamp_low[1]
port 54 nsew signal bidirectional
flabel metal3 s 324294 702300 326494 704800 0 FreeSans 1920 180 0 0 io_clamp_low[0]
port 53 nsew signal bidirectional
flabel metal3 s 173394 702300 175594 704800 0 FreeSans 1920 180 0 0 io_clamp_high[2]
port 52 nsew signal bidirectional
flabel metal3 s 225094 702300 227294 704800 0 FreeSans 1920 180 0 0 io_clamp_high[1]
port 51 nsew signal bidirectional
flabel metal3 s 326794 702300 328994 704800 0 FreeSans 1920 180 0 0 io_clamp_high[0]
port 50 nsew signal bidirectional
flabel metal5 s 217294 702300 222294 704800 0 FreeSans 1920 180 0 0 io_analog[5]
port 48 nsew signal bidirectional
flabel metal4 s 217294 702300 222294 704800 0 FreeSans 1920 180 0 0 io_analog[5]
port 48 nsew signal bidirectional
flabel metal3 s 217294 702300 222294 704800 0 FreeSans 1920 180 0 0 io_analog[5]
port 48 nsew signal bidirectional
flabel metal5 s 318994 702300 323994 704800 0 FreeSans 1920 180 0 0 io_analog[4]
port 47 nsew signal bidirectional
flabel metal4 s 318994 702300 323994 704800 0 FreeSans 1920 180 0 0 io_analog[4]
port 47 nsew signal bidirectional
flabel metal3 s 318994 702300 323994 704800 0 FreeSans 1920 180 0 0 io_analog[4]
port 47 nsew signal bidirectional
flabel metal3 s 16194 702300 21194 704800 0 FreeSans 1920 180 0 0 io_analog[9]
port 46 nsew signal bidirectional
flabel metal3 s 68194 702300 73194 704800 0 FreeSans 1920 180 0 0 io_analog[8]
port 45 nsew signal bidirectional
flabel metal3 s 120194 702300 125194 704800 0 FreeSans 1920 180 0 0 io_analog[7]
port 44 nsew signal bidirectional
flabel metal5 s 175894 702300 180894 704800 0 FreeSans 1920 180 0 0 io_analog[6]
port 43 nsew signal bidirectional
flabel metal5 s 227594 702300 232594 704800 0 FreeSans 1920 180 0 0 io_analog[5]
port 42 nsew signal bidirectional
flabel metal4 s 227594 702300 232594 704800 0 FreeSans 1920 180 0 0 io_analog[5]
port 42 nsew signal bidirectional
flabel metal3 s 227594 702300 232594 704800 0 FreeSans 1920 180 0 0 io_analog[5]
port 42 nsew signal bidirectional
flabel metal5 s 329294 702300 334294 704800 0 FreeSans 1920 180 0 0 io_analog[4]
port 41 nsew signal bidirectional
flabel metal4 s 329294 702300 334294 704800 0 FreeSans 1920 180 0 0 io_analog[4]
port 41 nsew signal bidirectional
flabel metal3 s 329294 702300 334294 704800 0 FreeSans 1920 180 0 0 io_analog[4]
port 41 nsew signal bidirectional
flabel metal3 s 413394 702300 418394 704800 0 FreeSans 1920 180 0 0 io_analog[3]
port 40 nsew signal bidirectional
flabel metal3 s 465394 702300 470394 704800 0 FreeSans 1920 180 0 0 io_analog[2]
port 39 nsew signal bidirectional
flabel metal3 s 566594 702300 571594 704800 0 FreeSans 1920 180 0 0 io_analog[1]
port 38 nsew signal bidirectional
flabel metal3 s 0 680242 1700 685242 0 FreeSans 1120 0 0 0 io_analog[10]
port 37 nsew signal bidirectional
flabel metal3 s 582300 677984 584800 682984 0 FreeSans 1120 0 0 0 io_analog[0]
port 36 nsew signal bidirectional
flabel metal3 s -800 423904 480 424016 0 FreeSans 1120 0 0 0 gpio_noesd[9]
port 35 nsew signal bidirectional
flabel metal3 s -800 467126 480 467238 0 FreeSans 1120 0 0 0 gpio_noesd[8]
port 34 nsew signal bidirectional
flabel metal3 s -800 510348 480 510460 0 FreeSans 1120 0 0 0 gpio_noesd[7]
port 33 nsew signal bidirectional
flabel metal3 s 583520 584744 584800 584856 0 FreeSans 1120 0 0 0 gpio_noesd[6]
port 32 nsew signal bidirectional
flabel metal3 s 583520 495322 584800 495434 0 FreeSans 1120 0 0 0 gpio_noesd[5]
port 31 nsew signal bidirectional
flabel metal3 s 583520 450900 584800 451012 0 FreeSans 1120 0 0 0 gpio_noesd[4]
port 30 nsew signal bidirectional
flabel metal3 s 583520 406478 584800 406590 0 FreeSans 1120 0 0 0 gpio_noesd[3]
port 29 nsew signal bidirectional
flabel metal3 s 583520 360056 584800 360168 0 FreeSans 1120 0 0 0 gpio_noesd[2]
port 28 nsew signal bidirectional
flabel metal3 s 583520 314834 584800 314946 0 FreeSans 1120 0 0 0 gpio_noesd[1]
port 27 nsew signal bidirectional
flabel metal3 s -800 15728 480 15840 0 FreeSans 1120 0 0 0 gpio_noesd[17]
port 26 nsew signal bidirectional
flabel metal3 s -800 37150 480 37262 0 FreeSans 1120 0 0 0 gpio_noesd[16]
port 25 nsew signal bidirectional
flabel metal3 s -800 80372 480 80484 0 FreeSans 1120 0 0 0 gpio_noesd[15]
port 24 nsew signal bidirectional
flabel metal3 s -800 123594 480 123706 0 FreeSans 1120 0 0 0 gpio_noesd[14]
port 23 nsew signal bidirectional
flabel metal3 s -800 251216 480 251328 0 FreeSans 1120 0 0 0 gpio_noesd[13]
port 22 nsew signal bidirectional
flabel metal3 s -800 294238 480 294350 0 FreeSans 1120 0 0 0 gpio_noesd[12]
port 21 nsew signal bidirectional
flabel metal3 s -800 337460 480 337572 0 FreeSans 1120 0 0 0 gpio_noesd[11]
port 20 nsew signal bidirectional
flabel metal3 s -800 380682 480 380794 0 FreeSans 1120 0 0 0 gpio_noesd[10]
port 19 nsew signal bidirectional
flabel metal3 s 583520 270412 584800 270524 0 FreeSans 1120 0 0 0 gpio_noesd[0]
port 18 nsew signal bidirectional
flabel metal3 s -800 425086 480 425198 0 FreeSans 1120 0 0 0 gpio_analog[9]
port 17 nsew signal bidirectional
flabel metal3 s -800 468308 480 468420 0 FreeSans 1120 0 0 0 gpio_analog[8]
port 16 nsew signal bidirectional
flabel metal3 s -800 511530 480 511642 0 FreeSans 1120 0 0 0 gpio_analog[7]
port 15 nsew signal bidirectional
flabel metal3 s 583520 583562 584800 583674 0 FreeSans 1120 0 0 0 gpio_analog[6]
port 14 nsew signal bidirectional
flabel metal3 s 583520 494140 584800 494252 0 FreeSans 1120 0 0 0 gpio_analog[5]
port 13 nsew signal bidirectional
flabel metal3 s 583520 449718 584800 449830 0 FreeSans 1120 0 0 0 gpio_analog[4]
port 12 nsew signal bidirectional
flabel metal3 s 583520 405296 584800 405408 0 FreeSans 1120 0 0 0 gpio_analog[3]
port 11 nsew signal bidirectional
flabel metal3 s 583520 358874 584800 358986 0 FreeSans 1120 0 0 0 gpio_analog[2]
port 10 nsew signal bidirectional
flabel metal3 s 583520 313652 584800 313764 0 FreeSans 1120 0 0 0 gpio_analog[1]
port 9 nsew signal bidirectional
flabel metal3 s -800 16910 480 17022 0 FreeSans 1120 0 0 0 gpio_analog[17]
port 8 nsew signal bidirectional
flabel metal3 s -800 38332 480 38444 0 FreeSans 1120 0 0 0 gpio_analog[16]
port 7 nsew signal bidirectional
flabel metal3 s -800 81554 480 81666 0 FreeSans 1120 0 0 0 gpio_analog[15]
port 6 nsew signal bidirectional
flabel metal3 s -800 124776 480 124888 0 FreeSans 1120 0 0 0 gpio_analog[14]
port 5 nsew signal bidirectional
flabel metal3 s -800 252398 480 252510 0 FreeSans 1120 0 0 0 gpio_analog[13]
port 4 nsew signal bidirectional
flabel metal3 s -800 295420 480 295532 0 FreeSans 1120 0 0 0 gpio_analog[12]
port 3 nsew signal bidirectional
flabel metal3 s -800 338642 480 338754 0 FreeSans 1120 0 0 0 gpio_analog[11]
port 2 nsew signal bidirectional
flabel metal3 s -800 381864 480 381976 0 FreeSans 1120 0 0 0 gpio_analog[10]
port 1 nsew signal bidirectional
flabel metal3 s 583520 269230 584800 269342 0 FreeSans 1120 0 0 0 gpio_analog[0]
port 0 nsew signal bidirectional
rlabel metal3 68306 691906 68306 691906 7 CLK
rlabel metal3 120364 698834 120364 698834 7 CLKBAR
rlabel metal3 413536 692644 413536 692644 7 Outn
rlabel metal3 469446 693308 469446 693308 3 Outp
rlabel metal4 552168 633194 552168 633194 5 VDD
rlabel metal5 524080 664482 524080 664482 3 GND
flabel metal5 s 165594 702300 170594 704800 0 FreeSans 1920 180 0 0 io_analog[6]
port 49 nsew signal bidirectional
flabel metal3 s 165596 702300 170596 704800 0 FreeSans 1920 180 0 0 io_analog[6]
port 49 nsew signal bidirectional
rlabel metal5 218258 702758 218258 702758 7 Vp
flabel metal3 s 175896 702300 180896 704800 0 FreeSans 1920 180 0 0 io_analog[6]
port 43 nsew signal bidirectional
rlabel metal5 166906 692944 166906 692944 7 Vn
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>
