magic
tech sky130A
timestamp 1651654828
<< end >>
